magic
tech scmos
timestamp 1732000943
<< nwell >>
rect -244 39 -220 91
rect -214 34 -190 89
rect -184 34 -160 89
rect -154 34 -130 89
rect -124 34 -100 89
rect -94 38 -70 90
rect -60 38 -36 90
rect -29 37 -5 89
rect 5 37 29 89
rect -214 -24 -190 28
rect -184 -24 -160 28
rect 43 -3 67 89
rect 73 -3 97 89
rect 103 37 127 89
rect 133 37 157 89
rect 163 37 187 89
rect 205 37 229 89
rect 235 37 259 89
rect 265 37 289 89
rect 311 -3 335 89
rect 370 37 394 89
rect 404 37 428 89
rect 453 -3 477 89
rect 483 -3 507 89
rect 513 37 537 89
rect 543 33 567 88
rect 573 33 597 88
rect 603 33 627 88
rect 633 33 657 88
rect 663 37 687 89
rect -89 -59 -65 -7
rect -55 -59 -31 -7
rect -24 -60 0 -8
rect 10 -60 34 -8
rect -241 -133 -217 -81
rect -211 -137 -187 -82
rect -181 -137 -157 -82
rect -151 -137 -127 -82
rect -121 -137 -97 -82
rect -211 -195 -187 -143
rect -181 -195 -157 -143
rect -88 -155 -64 -103
rect -54 -155 -30 -103
rect -23 -156 1 -104
rect 11 -156 35 -104
rect 43 -108 67 -16
rect 73 -108 97 -16
rect 103 -141 127 -89
rect 133 -141 157 -89
rect 163 -141 187 -89
rect 206 -141 230 -89
rect 236 -141 260 -89
rect 266 -141 290 -89
rect 311 -114 335 -22
rect 375 -60 399 -8
rect 409 -60 433 -8
rect 345 -113 369 -61
rect 376 -156 400 -104
rect 410 -156 434 -104
rect 453 -108 477 -16
rect 483 -108 507 -16
rect 543 -25 567 27
rect 573 -25 597 27
rect 513 -134 537 -82
rect 546 -138 570 -83
rect 576 -138 600 -83
rect 606 -138 630 -83
rect 636 -138 660 -83
rect 666 -134 690 -82
rect -243 -302 -219 -250
rect -213 -306 -189 -251
rect -183 -306 -159 -251
rect -153 -306 -129 -251
rect -123 -306 -99 -251
rect -83 -252 -59 -200
rect -49 -252 -25 -200
rect -18 -253 6 -201
rect 16 -253 40 -201
rect -213 -364 -189 -312
rect -183 -364 -159 -312
rect 47 -334 71 -242
rect 77 -334 101 -242
rect 311 -256 335 -164
rect 546 -196 570 -144
rect 576 -196 600 -144
rect 381 -253 405 -201
rect 415 -253 439 -201
rect 107 -319 131 -267
rect 137 -319 161 -267
rect 167 -319 191 -267
rect 202 -320 226 -268
rect 232 -320 256 -268
rect 262 -320 286 -268
rect -242 -471 -218 -419
rect -212 -475 -188 -420
rect -182 -475 -158 -420
rect -152 -475 -128 -420
rect -122 -475 -98 -420
rect 47 -439 71 -347
rect 77 -439 101 -347
rect 311 -367 335 -275
rect 345 -367 369 -315
rect 454 -334 478 -242
rect 484 -334 508 -242
rect 514 -303 538 -251
rect 544 -307 568 -252
rect 574 -307 598 -252
rect 604 -307 628 -252
rect 634 -307 658 -252
rect 664 -303 688 -251
rect -212 -533 -188 -481
rect -182 -533 -158 -481
rect 107 -497 131 -445
rect 137 -497 161 -445
rect 167 -497 191 -445
rect 203 -498 227 -446
rect 233 -498 257 -446
rect 263 -498 287 -446
rect 311 -509 335 -417
rect 454 -439 478 -347
rect 484 -439 508 -347
rect 544 -365 568 -313
rect 574 -365 598 -313
rect 514 -471 538 -419
rect 545 -476 569 -421
rect 575 -476 599 -421
rect 605 -476 629 -421
rect 635 -476 659 -421
rect 665 -472 689 -420
rect -237 -641 -213 -589
rect -207 -645 -183 -590
rect -177 -645 -153 -590
rect -147 -645 -123 -590
rect -117 -645 -93 -590
rect -207 -703 -183 -651
rect -177 -703 -153 -651
rect 52 -666 76 -574
rect 82 -666 106 -574
rect 311 -620 335 -528
rect 545 -534 569 -482
rect 575 -534 599 -482
rect 345 -620 369 -568
rect 455 -665 479 -573
rect 485 -665 509 -573
rect 515 -642 539 -590
rect 550 -646 574 -591
rect 580 -646 604 -591
rect 610 -646 634 -591
rect 640 -646 664 -591
rect 670 -642 694 -590
rect -234 -812 -210 -760
rect -204 -816 -180 -761
rect -174 -816 -150 -761
rect -144 -816 -120 -761
rect -114 -816 -90 -761
rect 52 -771 76 -679
rect 82 -771 106 -679
rect 311 -762 335 -670
rect 455 -770 479 -678
rect 485 -770 509 -678
rect 550 -704 574 -652
rect 580 -704 604 -652
rect -204 -874 -180 -822
rect -174 -874 -150 -822
rect 311 -873 335 -781
rect 345 -873 369 -821
rect -232 -983 -208 -931
rect -202 -987 -178 -932
rect -172 -987 -148 -932
rect -142 -987 -118 -932
rect -112 -987 -88 -932
rect -202 -1045 -178 -993
rect -172 -1045 -148 -993
rect 56 -999 80 -907
rect 86 -999 110 -907
rect 454 -996 478 -904
rect 484 -996 508 -904
rect -229 -1155 -205 -1103
rect 56 -1104 80 -1012
rect 86 -1104 110 -1012
rect 454 -1101 478 -1009
rect 484 -1101 508 -1009
rect -199 -1159 -175 -1104
rect -169 -1159 -145 -1104
rect -139 -1159 -115 -1104
rect -109 -1159 -85 -1104
rect -199 -1217 -175 -1165
rect -169 -1217 -145 -1165
<< ntransistor >>
rect -233 10 -231 30
rect -143 2 -141 22
rect -113 2 -111 22
rect -83 9 -81 29
rect -49 9 -47 29
rect -18 8 -16 28
rect 16 8 18 28
rect -143 -33 -141 -13
rect -113 -33 -111 -13
rect -203 -67 -201 -47
rect -173 -67 -171 -47
rect 114 -20 116 20
rect 174 8 176 28
rect 216 -20 218 20
rect 276 8 278 28
rect 381 8 383 28
rect 415 8 417 28
rect 524 8 526 28
rect -78 -88 -76 -68
rect -44 -88 -42 -68
rect -13 -89 -11 -69
rect 21 -89 23 -69
rect 114 -71 116 -31
rect 216 -71 218 -31
rect -230 -162 -228 -142
rect -140 -169 -138 -149
rect -110 -169 -108 -149
rect -77 -184 -75 -164
rect -43 -184 -41 -164
rect -140 -204 -138 -184
rect -110 -204 -108 -184
rect -12 -185 -10 -165
rect 22 -185 24 -165
rect 54 -169 56 -129
rect 84 -169 86 -129
rect 614 1 616 21
rect 644 1 646 21
rect 674 8 676 28
rect 386 -89 388 -69
rect 420 -89 422 -69
rect 614 -34 616 -14
rect 644 -34 646 -14
rect 554 -68 556 -48
rect 584 -68 586 -48
rect -200 -238 -198 -218
rect -170 -238 -168 -218
rect 54 -224 56 -184
rect 84 -224 86 -184
rect 114 -198 116 -158
rect 174 -170 176 -150
rect 217 -198 219 -158
rect 277 -170 279 -150
rect 322 -151 324 -131
rect 340 -151 342 -131
rect 356 -142 358 -122
rect -72 -281 -70 -261
rect -38 -281 -36 -261
rect -7 -282 -5 -262
rect 27 -282 29 -262
rect -232 -331 -230 -311
rect -142 -338 -140 -318
rect -112 -338 -110 -318
rect 114 -249 116 -209
rect 217 -249 219 -209
rect 387 -185 389 -165
rect 421 -185 423 -165
rect 464 -169 466 -129
rect 494 -169 496 -129
rect 524 -163 526 -143
rect 464 -224 466 -184
rect 494 -224 496 -184
rect 617 -170 619 -150
rect 647 -170 649 -150
rect 677 -163 679 -143
rect 617 -205 619 -185
rect 647 -205 649 -185
rect 557 -239 559 -219
rect 587 -239 589 -219
rect -142 -373 -140 -353
rect -112 -373 -110 -353
rect -202 -407 -200 -387
rect -172 -407 -170 -387
rect 118 -376 120 -336
rect 178 -348 180 -328
rect 213 -377 215 -337
rect 273 -349 275 -329
rect 392 -282 394 -262
rect 426 -282 428 -262
rect 525 -332 527 -312
rect 118 -427 120 -387
rect 213 -428 215 -388
rect 322 -404 324 -384
rect 340 -404 342 -384
rect 356 -396 358 -376
rect -231 -500 -229 -480
rect -141 -507 -139 -487
rect -111 -507 -109 -487
rect 58 -500 60 -460
rect 88 -500 90 -460
rect -141 -542 -139 -522
rect -111 -542 -109 -522
rect 58 -555 60 -515
rect 88 -555 90 -515
rect 118 -554 120 -514
rect 178 -526 180 -506
rect 615 -339 617 -319
rect 645 -339 647 -319
rect 675 -332 677 -312
rect 615 -374 617 -354
rect 645 -374 647 -354
rect 555 -408 557 -388
rect 585 -408 587 -388
rect 465 -500 467 -460
rect 495 -500 497 -460
rect 525 -500 527 -480
rect -201 -576 -199 -556
rect -171 -576 -169 -556
rect 214 -555 216 -515
rect 274 -527 276 -507
rect -226 -670 -224 -650
rect -136 -677 -134 -657
rect -106 -677 -104 -657
rect 118 -605 120 -565
rect 214 -606 216 -566
rect 465 -555 467 -515
rect 495 -555 497 -515
rect 616 -508 618 -488
rect 646 -508 648 -488
rect 676 -501 678 -481
rect 616 -543 618 -523
rect 646 -543 648 -523
rect 556 -577 558 -557
rect 586 -577 588 -557
rect 322 -657 324 -637
rect 340 -657 342 -637
rect 356 -649 358 -629
rect 526 -671 528 -651
rect -136 -712 -134 -692
rect -106 -712 -104 -692
rect -196 -746 -194 -726
rect -166 -746 -164 -726
rect 621 -678 623 -658
rect 651 -678 653 -658
rect 681 -671 683 -651
rect 621 -713 623 -693
rect 651 -713 653 -693
rect 561 -747 563 -727
rect 591 -747 593 -727
rect -223 -841 -221 -821
rect -133 -848 -131 -828
rect -103 -848 -101 -828
rect 63 -832 65 -792
rect 93 -832 95 -792
rect -133 -883 -131 -863
rect -103 -883 -101 -863
rect 63 -887 65 -847
rect 93 -887 95 -847
rect 466 -831 468 -791
rect 496 -831 498 -791
rect -193 -917 -191 -897
rect -163 -917 -161 -897
rect 322 -910 324 -890
rect 340 -910 342 -890
rect 356 -902 358 -882
rect 466 -886 468 -846
rect 496 -886 498 -846
rect -221 -1012 -219 -992
rect -131 -1019 -129 -999
rect -101 -1019 -99 -999
rect -131 -1054 -129 -1034
rect -101 -1054 -99 -1034
rect -191 -1088 -189 -1068
rect -161 -1088 -159 -1068
rect -218 -1184 -216 -1164
rect 67 -1165 69 -1125
rect 97 -1165 99 -1125
rect 465 -1162 467 -1122
rect 495 -1162 497 -1122
rect -128 -1191 -126 -1171
rect -98 -1191 -96 -1171
rect -128 -1226 -126 -1206
rect -98 -1226 -96 -1206
rect 67 -1220 69 -1180
rect 97 -1220 99 -1180
rect 465 -1217 467 -1177
rect 495 -1217 497 -1177
rect -188 -1260 -186 -1240
rect -158 -1260 -156 -1240
<< ptransistor >>
rect -233 45 -231 85
rect -203 43 -201 83
rect -173 43 -171 83
rect -143 43 -141 83
rect -113 43 -111 83
rect -83 44 -81 84
rect -49 44 -47 84
rect -18 43 -16 83
rect 16 43 18 83
rect -203 -18 -201 22
rect -173 -18 -171 22
rect 54 3 56 83
rect 84 3 86 83
rect 114 43 116 83
rect 144 43 146 83
rect 174 43 176 83
rect 216 43 218 83
rect 246 43 248 83
rect 276 43 278 83
rect -78 -53 -76 -13
rect -44 -53 -42 -13
rect -13 -54 -11 -14
rect 21 -54 23 -14
rect 322 3 324 83
rect 381 43 383 83
rect 415 43 417 83
rect 464 3 466 83
rect 494 3 496 83
rect 524 43 526 83
rect 554 42 556 82
rect 584 42 586 82
rect 614 42 616 82
rect 644 42 646 82
rect 674 43 676 83
rect -230 -127 -228 -87
rect -200 -128 -198 -88
rect -170 -128 -168 -88
rect -140 -128 -138 -88
rect -110 -128 -108 -88
rect 54 -102 56 -22
rect 84 -102 86 -22
rect -77 -149 -75 -109
rect -43 -149 -41 -109
rect -200 -189 -198 -149
rect -170 -189 -168 -149
rect -12 -150 -10 -110
rect 22 -150 24 -110
rect 114 -135 116 -95
rect 144 -135 146 -95
rect 174 -135 176 -95
rect 217 -135 219 -95
rect 247 -135 249 -95
rect 277 -135 279 -95
rect 322 -108 324 -28
rect 386 -54 388 -14
rect 420 -54 422 -14
rect 554 -19 556 21
rect 584 -19 586 21
rect 356 -107 358 -67
rect 464 -102 466 -22
rect 494 -102 496 -22
rect -72 -246 -70 -206
rect -38 -246 -36 -206
rect -232 -296 -230 -256
rect -202 -297 -200 -257
rect -172 -297 -170 -257
rect -142 -297 -140 -257
rect -112 -297 -110 -257
rect -7 -247 -5 -207
rect 27 -247 29 -207
rect 387 -150 389 -110
rect 421 -150 423 -110
rect 524 -128 526 -88
rect -202 -358 -200 -318
rect -172 -358 -170 -318
rect 58 -328 60 -248
rect 88 -328 90 -248
rect 322 -250 324 -170
rect 557 -129 559 -89
rect 587 -129 589 -89
rect 617 -129 619 -89
rect 647 -129 649 -89
rect 677 -128 679 -88
rect 392 -247 394 -207
rect 426 -247 428 -207
rect 557 -190 559 -150
rect 587 -190 589 -150
rect 118 -313 120 -273
rect 148 -313 150 -273
rect 178 -313 180 -273
rect 213 -314 215 -274
rect 243 -314 245 -274
rect 273 -314 275 -274
rect -231 -465 -229 -425
rect -201 -466 -199 -426
rect -171 -466 -169 -426
rect -141 -466 -139 -426
rect -111 -466 -109 -426
rect 58 -433 60 -353
rect 88 -433 90 -353
rect 322 -361 324 -281
rect 356 -361 358 -321
rect 465 -328 467 -248
rect 495 -328 497 -248
rect 525 -297 527 -257
rect 555 -298 557 -258
rect 585 -298 587 -258
rect 615 -298 617 -258
rect 645 -298 647 -258
rect 675 -297 677 -257
rect -201 -527 -199 -487
rect -171 -527 -169 -487
rect 118 -491 120 -451
rect 148 -491 150 -451
rect 178 -491 180 -451
rect 214 -492 216 -452
rect 244 -492 246 -452
rect 274 -492 276 -452
rect 322 -503 324 -423
rect 465 -433 467 -353
rect 495 -433 497 -353
rect 555 -359 557 -319
rect 585 -359 587 -319
rect 525 -465 527 -425
rect 556 -467 558 -427
rect 586 -467 588 -427
rect 616 -467 618 -427
rect 646 -467 648 -427
rect 676 -466 678 -426
rect -226 -635 -224 -595
rect -196 -636 -194 -596
rect -166 -636 -164 -596
rect -136 -636 -134 -596
rect -106 -636 -104 -596
rect -196 -697 -194 -657
rect -166 -697 -164 -657
rect 63 -660 65 -580
rect 93 -660 95 -580
rect 322 -614 324 -534
rect 556 -528 558 -488
rect 586 -528 588 -488
rect 356 -614 358 -574
rect 466 -659 468 -579
rect 496 -659 498 -579
rect 526 -636 528 -596
rect 561 -637 563 -597
rect 591 -637 593 -597
rect 621 -637 623 -597
rect 651 -637 653 -597
rect 681 -636 683 -596
rect -223 -806 -221 -766
rect 63 -765 65 -685
rect 93 -765 95 -685
rect 322 -756 324 -676
rect -193 -807 -191 -767
rect -163 -807 -161 -767
rect -133 -807 -131 -767
rect -103 -807 -101 -767
rect 466 -764 468 -684
rect 496 -764 498 -684
rect 561 -698 563 -658
rect 591 -698 593 -658
rect -193 -868 -191 -828
rect -163 -868 -161 -828
rect 322 -867 324 -787
rect 356 -867 358 -827
rect -221 -977 -219 -937
rect -191 -978 -189 -938
rect -161 -978 -159 -938
rect -131 -978 -129 -938
rect -101 -978 -99 -938
rect 67 -993 69 -913
rect 97 -993 99 -913
rect 465 -990 467 -910
rect 495 -990 497 -910
rect -191 -1039 -189 -999
rect -161 -1039 -159 -999
rect 67 -1098 69 -1018
rect 97 -1098 99 -1018
rect 465 -1095 467 -1015
rect 495 -1095 497 -1015
rect -218 -1149 -216 -1109
rect -188 -1150 -186 -1110
rect -158 -1150 -156 -1110
rect -128 -1150 -126 -1110
rect -98 -1150 -96 -1110
rect -188 -1211 -186 -1171
rect -158 -1211 -156 -1171
<< ndiffusion >>
rect -234 10 -233 30
rect -231 10 -230 30
rect -144 2 -143 22
rect -141 2 -140 22
rect -114 2 -113 22
rect -111 2 -110 22
rect -84 9 -83 29
rect -81 9 -80 29
rect -50 9 -49 29
rect -47 9 -46 29
rect -19 8 -18 28
rect -16 8 -15 28
rect 15 8 16 28
rect 18 8 19 28
rect -144 -33 -143 -13
rect -141 -33 -140 -13
rect -114 -33 -113 -13
rect -111 -33 -110 -13
rect -204 -67 -203 -47
rect -201 -67 -200 -47
rect -174 -67 -173 -47
rect -171 -67 -170 -47
rect 113 -20 114 20
rect 116 -20 117 20
rect 173 8 174 28
rect 176 8 177 28
rect 215 -20 216 20
rect 218 -20 219 20
rect 275 8 276 28
rect 278 8 279 28
rect 380 8 381 28
rect 383 8 384 28
rect 414 8 415 28
rect 417 8 418 28
rect 523 8 524 28
rect 526 8 527 28
rect -79 -88 -78 -68
rect -76 -88 -75 -68
rect -45 -88 -44 -68
rect -42 -88 -41 -68
rect -14 -89 -13 -69
rect -11 -89 -10 -69
rect 20 -89 21 -69
rect 23 -89 24 -69
rect 113 -71 114 -31
rect 116 -71 117 -31
rect 215 -71 216 -31
rect 218 -71 219 -31
rect -231 -162 -230 -142
rect -228 -162 -227 -142
rect -141 -169 -140 -149
rect -138 -169 -137 -149
rect -111 -169 -110 -149
rect -108 -169 -107 -149
rect -78 -184 -77 -164
rect -75 -184 -74 -164
rect -44 -184 -43 -164
rect -41 -184 -40 -164
rect -141 -204 -140 -184
rect -138 -204 -137 -184
rect -111 -204 -110 -184
rect -108 -204 -107 -184
rect -13 -185 -12 -165
rect -10 -185 -9 -165
rect 21 -185 22 -165
rect 24 -185 25 -165
rect 53 -169 54 -129
rect 56 -169 57 -129
rect 83 -169 84 -129
rect 86 -169 87 -129
rect 613 1 614 21
rect 616 1 617 21
rect 643 1 644 21
rect 646 1 647 21
rect 673 8 674 28
rect 676 8 677 28
rect 385 -89 386 -69
rect 388 -89 389 -69
rect 419 -89 420 -69
rect 422 -89 423 -69
rect 613 -34 614 -14
rect 616 -34 617 -14
rect 643 -34 644 -14
rect 646 -34 647 -14
rect 553 -68 554 -48
rect 556 -68 557 -48
rect 583 -68 584 -48
rect 586 -68 587 -48
rect -201 -238 -200 -218
rect -198 -238 -197 -218
rect -171 -238 -170 -218
rect -168 -238 -167 -218
rect 53 -224 54 -184
rect 56 -224 57 -184
rect 83 -224 84 -184
rect 86 -224 87 -184
rect 113 -198 114 -158
rect 116 -198 117 -158
rect 173 -170 174 -150
rect 176 -170 177 -150
rect 216 -198 217 -158
rect 219 -198 220 -158
rect 276 -170 277 -150
rect 279 -170 280 -150
rect 321 -151 322 -131
rect 324 -151 325 -131
rect 339 -151 340 -131
rect 342 -151 343 -131
rect 355 -142 356 -122
rect 358 -142 359 -122
rect -73 -281 -72 -261
rect -70 -281 -69 -261
rect -39 -281 -38 -261
rect -36 -281 -35 -261
rect -8 -282 -7 -262
rect -5 -282 -4 -262
rect 26 -282 27 -262
rect 29 -282 30 -262
rect -233 -331 -232 -311
rect -230 -331 -229 -311
rect -143 -338 -142 -318
rect -140 -338 -139 -318
rect -113 -338 -112 -318
rect -110 -338 -109 -318
rect 113 -249 114 -209
rect 116 -249 117 -209
rect 216 -249 217 -209
rect 219 -249 220 -209
rect 386 -185 387 -165
rect 389 -185 390 -165
rect 420 -185 421 -165
rect 423 -185 424 -165
rect 463 -169 464 -129
rect 466 -169 467 -129
rect 493 -169 494 -129
rect 496 -169 497 -129
rect 523 -163 524 -143
rect 526 -163 527 -143
rect 463 -224 464 -184
rect 466 -224 467 -184
rect 493 -224 494 -184
rect 496 -224 497 -184
rect 616 -170 617 -150
rect 619 -170 620 -150
rect 646 -170 647 -150
rect 649 -170 650 -150
rect 676 -163 677 -143
rect 679 -163 680 -143
rect 616 -205 617 -185
rect 619 -205 620 -185
rect 646 -205 647 -185
rect 649 -205 650 -185
rect 556 -239 557 -219
rect 559 -239 560 -219
rect 586 -239 587 -219
rect 589 -239 590 -219
rect -143 -373 -142 -353
rect -140 -373 -139 -353
rect -113 -373 -112 -353
rect -110 -373 -109 -353
rect -203 -407 -202 -387
rect -200 -407 -199 -387
rect -173 -407 -172 -387
rect -170 -407 -169 -387
rect 117 -376 118 -336
rect 120 -376 121 -336
rect 177 -348 178 -328
rect 180 -348 181 -328
rect 212 -377 213 -337
rect 215 -377 216 -337
rect 272 -349 273 -329
rect 275 -349 276 -329
rect 391 -282 392 -262
rect 394 -282 395 -262
rect 425 -282 426 -262
rect 428 -282 429 -262
rect 524 -332 525 -312
rect 527 -332 528 -312
rect 117 -427 118 -387
rect 120 -427 121 -387
rect 212 -428 213 -388
rect 215 -428 216 -388
rect 321 -404 322 -384
rect 324 -404 325 -384
rect 339 -404 340 -384
rect 342 -404 343 -384
rect 355 -396 356 -376
rect 358 -396 359 -376
rect -232 -500 -231 -480
rect -229 -500 -228 -480
rect -142 -507 -141 -487
rect -139 -507 -138 -487
rect -112 -507 -111 -487
rect -109 -507 -108 -487
rect 57 -500 58 -460
rect 60 -500 61 -460
rect 87 -500 88 -460
rect 90 -500 91 -460
rect -142 -542 -141 -522
rect -139 -542 -138 -522
rect -112 -542 -111 -522
rect -109 -542 -108 -522
rect 57 -555 58 -515
rect 60 -555 61 -515
rect 87 -555 88 -515
rect 90 -555 91 -515
rect 117 -554 118 -514
rect 120 -554 121 -514
rect 177 -526 178 -506
rect 180 -526 181 -506
rect 614 -339 615 -319
rect 617 -339 618 -319
rect 644 -339 645 -319
rect 647 -339 648 -319
rect 674 -332 675 -312
rect 677 -332 678 -312
rect 614 -374 615 -354
rect 617 -374 618 -354
rect 644 -374 645 -354
rect 647 -374 648 -354
rect 554 -408 555 -388
rect 557 -408 558 -388
rect 584 -408 585 -388
rect 587 -408 588 -388
rect 464 -500 465 -460
rect 467 -500 468 -460
rect 494 -500 495 -460
rect 497 -500 498 -460
rect 524 -500 525 -480
rect 527 -500 528 -480
rect -202 -576 -201 -556
rect -199 -576 -198 -556
rect -172 -576 -171 -556
rect -169 -576 -168 -556
rect 213 -555 214 -515
rect 216 -555 217 -515
rect 273 -527 274 -507
rect 276 -527 277 -507
rect -227 -670 -226 -650
rect -224 -670 -223 -650
rect -137 -677 -136 -657
rect -134 -677 -133 -657
rect -107 -677 -106 -657
rect -104 -677 -103 -657
rect 117 -605 118 -565
rect 120 -605 121 -565
rect 213 -606 214 -566
rect 216 -606 217 -566
rect 464 -555 465 -515
rect 467 -555 468 -515
rect 494 -555 495 -515
rect 497 -555 498 -515
rect 615 -508 616 -488
rect 618 -508 619 -488
rect 645 -508 646 -488
rect 648 -508 649 -488
rect 675 -501 676 -481
rect 678 -501 679 -481
rect 615 -543 616 -523
rect 618 -543 619 -523
rect 645 -543 646 -523
rect 648 -543 649 -523
rect 555 -577 556 -557
rect 558 -577 559 -557
rect 585 -577 586 -557
rect 588 -577 589 -557
rect 321 -657 322 -637
rect 324 -657 325 -637
rect 339 -657 340 -637
rect 342 -657 343 -637
rect 355 -649 356 -629
rect 358 -649 359 -629
rect 525 -671 526 -651
rect 528 -671 529 -651
rect -137 -712 -136 -692
rect -134 -712 -133 -692
rect -107 -712 -106 -692
rect -104 -712 -103 -692
rect -197 -746 -196 -726
rect -194 -746 -193 -726
rect -167 -746 -166 -726
rect -164 -746 -163 -726
rect 620 -678 621 -658
rect 623 -678 624 -658
rect 650 -678 651 -658
rect 653 -678 654 -658
rect 680 -671 681 -651
rect 683 -671 684 -651
rect 620 -713 621 -693
rect 623 -713 624 -693
rect 650 -713 651 -693
rect 653 -713 654 -693
rect 560 -747 561 -727
rect 563 -747 564 -727
rect 590 -747 591 -727
rect 593 -747 594 -727
rect -224 -841 -223 -821
rect -221 -841 -220 -821
rect -134 -848 -133 -828
rect -131 -848 -130 -828
rect -104 -848 -103 -828
rect -101 -848 -100 -828
rect 62 -832 63 -792
rect 65 -832 66 -792
rect 92 -832 93 -792
rect 95 -832 96 -792
rect -134 -883 -133 -863
rect -131 -883 -130 -863
rect -104 -883 -103 -863
rect -101 -883 -100 -863
rect 62 -887 63 -847
rect 65 -887 66 -847
rect 92 -887 93 -847
rect 95 -887 96 -847
rect 465 -831 466 -791
rect 468 -831 469 -791
rect 495 -831 496 -791
rect 498 -831 499 -791
rect -194 -917 -193 -897
rect -191 -917 -190 -897
rect -164 -917 -163 -897
rect -161 -917 -160 -897
rect 321 -910 322 -890
rect 324 -910 325 -890
rect 339 -910 340 -890
rect 342 -910 343 -890
rect 355 -902 356 -882
rect 358 -902 359 -882
rect 465 -886 466 -846
rect 468 -886 469 -846
rect 495 -886 496 -846
rect 498 -886 499 -846
rect -222 -1012 -221 -992
rect -219 -1012 -218 -992
rect -132 -1019 -131 -999
rect -129 -1019 -128 -999
rect -102 -1019 -101 -999
rect -99 -1019 -98 -999
rect -132 -1054 -131 -1034
rect -129 -1054 -128 -1034
rect -102 -1054 -101 -1034
rect -99 -1054 -98 -1034
rect -192 -1088 -191 -1068
rect -189 -1088 -188 -1068
rect -162 -1088 -161 -1068
rect -159 -1088 -158 -1068
rect -219 -1184 -218 -1164
rect -216 -1184 -215 -1164
rect 66 -1165 67 -1125
rect 69 -1165 70 -1125
rect 96 -1165 97 -1125
rect 99 -1165 100 -1125
rect 464 -1162 465 -1122
rect 467 -1162 468 -1122
rect 494 -1162 495 -1122
rect 497 -1162 498 -1122
rect -129 -1191 -128 -1171
rect -126 -1191 -125 -1171
rect -99 -1191 -98 -1171
rect -96 -1191 -95 -1171
rect -129 -1226 -128 -1206
rect -126 -1226 -125 -1206
rect -99 -1226 -98 -1206
rect -96 -1226 -95 -1206
rect 66 -1220 67 -1180
rect 69 -1220 70 -1180
rect 96 -1220 97 -1180
rect 99 -1220 100 -1180
rect 464 -1217 465 -1177
rect 467 -1217 468 -1177
rect 494 -1217 495 -1177
rect 497 -1217 498 -1177
rect -189 -1260 -188 -1240
rect -186 -1260 -185 -1240
rect -159 -1260 -158 -1240
rect -156 -1260 -155 -1240
<< pdiffusion >>
rect -234 45 -233 85
rect -231 45 -230 85
rect -204 43 -203 83
rect -201 43 -200 83
rect -174 43 -173 83
rect -171 43 -170 83
rect -144 43 -143 83
rect -141 43 -140 83
rect -114 43 -113 83
rect -111 43 -110 83
rect -84 44 -83 84
rect -81 44 -80 84
rect -50 44 -49 84
rect -47 44 -46 84
rect -19 43 -18 83
rect -16 43 -15 83
rect 15 43 16 83
rect 18 43 19 83
rect -204 -18 -203 22
rect -201 -18 -200 22
rect -174 -18 -173 22
rect -171 -18 -170 22
rect 53 3 54 83
rect 56 3 57 83
rect 83 3 84 83
rect 86 3 87 83
rect 113 43 114 83
rect 116 43 117 83
rect 143 43 144 83
rect 146 43 147 83
rect 173 43 174 83
rect 176 43 177 83
rect 215 43 216 83
rect 218 43 219 83
rect 245 43 246 83
rect 248 43 249 83
rect 275 43 276 83
rect 278 43 279 83
rect -79 -53 -78 -13
rect -76 -53 -75 -13
rect -45 -53 -44 -13
rect -42 -53 -41 -13
rect -14 -54 -13 -14
rect -11 -54 -10 -14
rect 20 -54 21 -14
rect 23 -54 24 -14
rect 321 3 322 83
rect 324 3 325 83
rect 380 43 381 83
rect 383 43 384 83
rect 414 43 415 83
rect 417 43 418 83
rect 463 3 464 83
rect 466 3 467 83
rect 493 3 494 83
rect 496 3 497 83
rect 523 43 524 83
rect 526 43 527 83
rect 553 42 554 82
rect 556 42 557 82
rect 583 42 584 82
rect 586 42 587 82
rect 613 42 614 82
rect 616 42 617 82
rect 643 42 644 82
rect 646 42 647 82
rect 673 43 674 83
rect 676 43 677 83
rect -231 -127 -230 -87
rect -228 -127 -227 -87
rect -201 -128 -200 -88
rect -198 -128 -197 -88
rect -171 -128 -170 -88
rect -168 -128 -167 -88
rect -141 -128 -140 -88
rect -138 -128 -137 -88
rect -111 -128 -110 -88
rect -108 -128 -107 -88
rect 53 -102 54 -22
rect 56 -102 57 -22
rect 83 -102 84 -22
rect 86 -102 87 -22
rect -78 -149 -77 -109
rect -75 -149 -74 -109
rect -44 -149 -43 -109
rect -41 -149 -40 -109
rect -201 -189 -200 -149
rect -198 -189 -197 -149
rect -171 -189 -170 -149
rect -168 -189 -167 -149
rect -13 -150 -12 -110
rect -10 -150 -9 -110
rect 21 -150 22 -110
rect 24 -150 25 -110
rect 113 -135 114 -95
rect 116 -135 117 -95
rect 143 -135 144 -95
rect 146 -135 147 -95
rect 173 -135 174 -95
rect 176 -135 177 -95
rect 216 -135 217 -95
rect 219 -135 220 -95
rect 246 -135 247 -95
rect 249 -135 250 -95
rect 276 -135 277 -95
rect 279 -135 280 -95
rect 321 -108 322 -28
rect 324 -108 325 -28
rect 385 -54 386 -14
rect 388 -54 389 -14
rect 419 -54 420 -14
rect 422 -54 423 -14
rect 553 -19 554 21
rect 556 -19 557 21
rect 583 -19 584 21
rect 586 -19 587 21
rect 355 -107 356 -67
rect 358 -107 359 -67
rect 463 -102 464 -22
rect 466 -102 467 -22
rect 493 -102 494 -22
rect 496 -102 497 -22
rect -73 -246 -72 -206
rect -70 -246 -69 -206
rect -39 -246 -38 -206
rect -36 -246 -35 -206
rect -233 -296 -232 -256
rect -230 -296 -229 -256
rect -203 -297 -202 -257
rect -200 -297 -199 -257
rect -173 -297 -172 -257
rect -170 -297 -169 -257
rect -143 -297 -142 -257
rect -140 -297 -139 -257
rect -113 -297 -112 -257
rect -110 -297 -109 -257
rect -8 -247 -7 -207
rect -5 -247 -4 -207
rect 26 -247 27 -207
rect 29 -247 30 -207
rect 386 -150 387 -110
rect 389 -150 390 -110
rect 420 -150 421 -110
rect 423 -150 424 -110
rect 523 -128 524 -88
rect 526 -128 527 -88
rect -203 -358 -202 -318
rect -200 -358 -199 -318
rect -173 -358 -172 -318
rect -170 -358 -169 -318
rect 57 -328 58 -248
rect 60 -328 61 -248
rect 87 -328 88 -248
rect 90 -328 91 -248
rect 321 -250 322 -170
rect 324 -250 325 -170
rect 556 -129 557 -89
rect 559 -129 560 -89
rect 586 -129 587 -89
rect 589 -129 590 -89
rect 616 -129 617 -89
rect 619 -129 620 -89
rect 646 -129 647 -89
rect 649 -129 650 -89
rect 676 -128 677 -88
rect 679 -128 680 -88
rect 391 -247 392 -207
rect 394 -247 395 -207
rect 425 -247 426 -207
rect 428 -247 429 -207
rect 556 -190 557 -150
rect 559 -190 560 -150
rect 586 -190 587 -150
rect 589 -190 590 -150
rect 117 -313 118 -273
rect 120 -313 121 -273
rect 147 -313 148 -273
rect 150 -313 151 -273
rect 177 -313 178 -273
rect 180 -313 181 -273
rect 212 -314 213 -274
rect 215 -314 216 -274
rect 242 -314 243 -274
rect 245 -314 246 -274
rect 272 -314 273 -274
rect 275 -314 276 -274
rect -232 -465 -231 -425
rect -229 -465 -228 -425
rect -202 -466 -201 -426
rect -199 -466 -198 -426
rect -172 -466 -171 -426
rect -169 -466 -168 -426
rect -142 -466 -141 -426
rect -139 -466 -138 -426
rect -112 -466 -111 -426
rect -109 -466 -108 -426
rect 57 -433 58 -353
rect 60 -433 61 -353
rect 87 -433 88 -353
rect 90 -433 91 -353
rect 321 -361 322 -281
rect 324 -361 325 -281
rect 355 -361 356 -321
rect 358 -361 359 -321
rect 464 -328 465 -248
rect 467 -328 468 -248
rect 494 -328 495 -248
rect 497 -328 498 -248
rect 524 -297 525 -257
rect 527 -297 528 -257
rect 554 -298 555 -258
rect 557 -298 558 -258
rect 584 -298 585 -258
rect 587 -298 588 -258
rect 614 -298 615 -258
rect 617 -298 618 -258
rect 644 -298 645 -258
rect 647 -298 648 -258
rect 674 -297 675 -257
rect 677 -297 678 -257
rect -202 -527 -201 -487
rect -199 -527 -198 -487
rect -172 -527 -171 -487
rect -169 -527 -168 -487
rect 117 -491 118 -451
rect 120 -491 121 -451
rect 147 -491 148 -451
rect 150 -491 151 -451
rect 177 -491 178 -451
rect 180 -491 181 -451
rect 213 -492 214 -452
rect 216 -492 217 -452
rect 243 -492 244 -452
rect 246 -492 247 -452
rect 273 -492 274 -452
rect 276 -492 277 -452
rect 321 -503 322 -423
rect 324 -503 325 -423
rect 464 -433 465 -353
rect 467 -433 468 -353
rect 494 -433 495 -353
rect 497 -433 498 -353
rect 554 -359 555 -319
rect 557 -359 558 -319
rect 584 -359 585 -319
rect 587 -359 588 -319
rect 524 -465 525 -425
rect 527 -465 528 -425
rect 555 -467 556 -427
rect 558 -467 559 -427
rect 585 -467 586 -427
rect 588 -467 589 -427
rect 615 -467 616 -427
rect 618 -467 619 -427
rect 645 -467 646 -427
rect 648 -467 649 -427
rect 675 -466 676 -426
rect 678 -466 679 -426
rect -227 -635 -226 -595
rect -224 -635 -223 -595
rect -197 -636 -196 -596
rect -194 -636 -193 -596
rect -167 -636 -166 -596
rect -164 -636 -163 -596
rect -137 -636 -136 -596
rect -134 -636 -133 -596
rect -107 -636 -106 -596
rect -104 -636 -103 -596
rect -197 -697 -196 -657
rect -194 -697 -193 -657
rect -167 -697 -166 -657
rect -164 -697 -163 -657
rect 62 -660 63 -580
rect 65 -660 66 -580
rect 92 -660 93 -580
rect 95 -660 96 -580
rect 321 -614 322 -534
rect 324 -614 325 -534
rect 555 -528 556 -488
rect 558 -528 559 -488
rect 585 -528 586 -488
rect 588 -528 589 -488
rect 355 -614 356 -574
rect 358 -614 359 -574
rect 465 -659 466 -579
rect 468 -659 469 -579
rect 495 -659 496 -579
rect 498 -659 499 -579
rect 525 -636 526 -596
rect 528 -636 529 -596
rect 560 -637 561 -597
rect 563 -637 564 -597
rect 590 -637 591 -597
rect 593 -637 594 -597
rect 620 -637 621 -597
rect 623 -637 624 -597
rect 650 -637 651 -597
rect 653 -637 654 -597
rect 680 -636 681 -596
rect 683 -636 684 -596
rect -224 -806 -223 -766
rect -221 -806 -220 -766
rect 62 -765 63 -685
rect 65 -765 66 -685
rect 92 -765 93 -685
rect 95 -765 96 -685
rect 321 -756 322 -676
rect 324 -756 325 -676
rect -194 -807 -193 -767
rect -191 -807 -190 -767
rect -164 -807 -163 -767
rect -161 -807 -160 -767
rect -134 -807 -133 -767
rect -131 -807 -130 -767
rect -104 -807 -103 -767
rect -101 -807 -100 -767
rect 465 -764 466 -684
rect 468 -764 469 -684
rect 495 -764 496 -684
rect 498 -764 499 -684
rect 560 -698 561 -658
rect 563 -698 564 -658
rect 590 -698 591 -658
rect 593 -698 594 -658
rect -194 -868 -193 -828
rect -191 -868 -190 -828
rect -164 -868 -163 -828
rect -161 -868 -160 -828
rect 321 -867 322 -787
rect 324 -867 325 -787
rect 355 -867 356 -827
rect 358 -867 359 -827
rect -222 -977 -221 -937
rect -219 -977 -218 -937
rect -192 -978 -191 -938
rect -189 -978 -188 -938
rect -162 -978 -161 -938
rect -159 -978 -158 -938
rect -132 -978 -131 -938
rect -129 -978 -128 -938
rect -102 -978 -101 -938
rect -99 -978 -98 -938
rect 66 -993 67 -913
rect 69 -993 70 -913
rect 96 -993 97 -913
rect 99 -993 100 -913
rect 464 -990 465 -910
rect 467 -990 468 -910
rect 494 -990 495 -910
rect 497 -990 498 -910
rect -192 -1039 -191 -999
rect -189 -1039 -188 -999
rect -162 -1039 -161 -999
rect -159 -1039 -158 -999
rect 66 -1098 67 -1018
rect 69 -1098 70 -1018
rect 96 -1098 97 -1018
rect 99 -1098 100 -1018
rect 464 -1095 465 -1015
rect 467 -1095 468 -1015
rect 494 -1095 495 -1015
rect 497 -1095 498 -1015
rect -219 -1149 -218 -1109
rect -216 -1149 -215 -1109
rect -189 -1150 -188 -1110
rect -186 -1150 -185 -1110
rect -159 -1150 -158 -1110
rect -156 -1150 -155 -1110
rect -129 -1150 -128 -1110
rect -126 -1150 -125 -1110
rect -99 -1150 -98 -1110
rect -96 -1150 -95 -1110
rect -189 -1211 -188 -1171
rect -186 -1211 -185 -1171
rect -159 -1211 -158 -1171
rect -156 -1211 -155 -1171
<< ndcontact >>
rect -238 10 -234 30
rect -230 10 -226 30
rect -148 2 -144 22
rect -140 2 -136 22
rect -118 2 -114 22
rect -110 2 -106 22
rect -88 9 -84 29
rect -80 9 -76 29
rect -54 9 -50 29
rect -46 9 -42 29
rect -23 8 -19 28
rect -15 8 -11 28
rect 11 8 15 28
rect 19 8 23 28
rect -148 -33 -144 -13
rect -140 -33 -136 -13
rect -118 -33 -114 -13
rect -110 -33 -106 -13
rect -208 -67 -204 -47
rect -200 -67 -196 -47
rect -178 -67 -174 -47
rect -170 -67 -166 -47
rect 109 -20 113 20
rect 117 -20 121 20
rect 169 8 173 28
rect 177 8 181 28
rect 211 -20 215 20
rect 219 -20 223 20
rect 271 8 275 28
rect 279 8 283 28
rect 376 8 380 28
rect 384 8 388 28
rect 410 8 414 28
rect 418 8 422 28
rect 519 8 523 28
rect 527 8 531 28
rect -83 -88 -79 -68
rect -75 -88 -71 -68
rect -49 -88 -45 -68
rect -41 -88 -37 -68
rect -18 -89 -14 -69
rect -10 -89 -6 -69
rect 16 -89 20 -69
rect 24 -89 28 -69
rect 109 -71 113 -31
rect 117 -71 121 -31
rect 211 -71 215 -31
rect 219 -71 223 -31
rect -235 -162 -231 -142
rect -227 -162 -223 -142
rect -145 -169 -141 -149
rect -137 -169 -133 -149
rect -115 -169 -111 -149
rect -107 -169 -103 -149
rect -82 -184 -78 -164
rect -74 -184 -70 -164
rect -48 -184 -44 -164
rect -40 -184 -36 -164
rect -145 -204 -141 -184
rect -137 -204 -133 -184
rect -115 -204 -111 -184
rect -107 -204 -103 -184
rect -17 -185 -13 -165
rect -9 -185 -5 -165
rect 17 -185 21 -165
rect 25 -185 29 -165
rect 49 -169 53 -129
rect 57 -169 61 -129
rect 79 -169 83 -129
rect 87 -169 91 -129
rect 609 1 613 21
rect 617 1 621 21
rect 639 1 643 21
rect 647 1 651 21
rect 669 8 673 28
rect 677 8 681 28
rect 381 -89 385 -69
rect 389 -89 393 -69
rect 415 -89 419 -69
rect 423 -89 427 -69
rect 609 -34 613 -14
rect 617 -34 621 -14
rect 639 -34 643 -14
rect 647 -34 651 -14
rect 549 -68 553 -48
rect 557 -68 561 -48
rect 579 -68 583 -48
rect 587 -68 591 -48
rect -205 -238 -201 -218
rect -197 -238 -193 -218
rect -175 -238 -171 -218
rect -167 -238 -163 -218
rect 49 -224 53 -184
rect 57 -224 61 -184
rect 79 -224 83 -184
rect 87 -224 91 -184
rect 109 -198 113 -158
rect 117 -198 121 -158
rect 169 -170 173 -150
rect 177 -170 181 -150
rect 212 -198 216 -158
rect 220 -198 224 -158
rect 272 -170 276 -150
rect 280 -170 284 -150
rect 317 -151 321 -131
rect 325 -151 329 -131
rect 335 -151 339 -131
rect 343 -151 347 -131
rect 351 -142 355 -122
rect 359 -142 363 -122
rect -77 -281 -73 -261
rect -69 -281 -65 -261
rect -43 -281 -39 -261
rect -35 -281 -31 -261
rect -12 -282 -8 -262
rect -4 -282 0 -262
rect 22 -282 26 -262
rect 30 -282 34 -262
rect -237 -331 -233 -311
rect -229 -331 -225 -311
rect -147 -338 -143 -318
rect -139 -338 -135 -318
rect -117 -338 -113 -318
rect -109 -338 -105 -318
rect 109 -249 113 -209
rect 117 -249 121 -209
rect 212 -249 216 -209
rect 220 -249 224 -209
rect 382 -185 386 -165
rect 390 -185 394 -165
rect 416 -185 420 -165
rect 424 -185 428 -165
rect 459 -169 463 -129
rect 467 -169 471 -129
rect 489 -169 493 -129
rect 497 -169 501 -129
rect 519 -163 523 -143
rect 527 -163 531 -143
rect 459 -224 463 -184
rect 467 -224 471 -184
rect 489 -224 493 -184
rect 497 -224 501 -184
rect 612 -170 616 -150
rect 620 -170 624 -150
rect 642 -170 646 -150
rect 650 -170 654 -150
rect 672 -163 676 -143
rect 680 -163 684 -143
rect 612 -205 616 -185
rect 620 -205 624 -185
rect 642 -205 646 -185
rect 650 -205 654 -185
rect 552 -239 556 -219
rect 560 -239 564 -219
rect 582 -239 586 -219
rect 590 -239 594 -219
rect -147 -373 -143 -353
rect -139 -373 -135 -353
rect -117 -373 -113 -353
rect -109 -373 -105 -353
rect -207 -407 -203 -387
rect -199 -407 -195 -387
rect -177 -407 -173 -387
rect -169 -407 -165 -387
rect 113 -376 117 -336
rect 121 -376 125 -336
rect 173 -348 177 -328
rect 181 -348 185 -328
rect 208 -377 212 -337
rect 216 -377 220 -337
rect 268 -349 272 -329
rect 276 -349 280 -329
rect 387 -282 391 -262
rect 395 -282 399 -262
rect 421 -282 425 -262
rect 429 -282 433 -262
rect 520 -332 524 -312
rect 528 -332 532 -312
rect 113 -427 117 -387
rect 121 -427 125 -387
rect 208 -428 212 -388
rect 216 -428 220 -388
rect 317 -404 321 -384
rect 325 -404 329 -384
rect 335 -404 339 -384
rect 343 -404 347 -384
rect 351 -396 355 -376
rect 359 -396 363 -376
rect -236 -500 -232 -480
rect -228 -500 -224 -480
rect -146 -507 -142 -487
rect -138 -507 -134 -487
rect -116 -507 -112 -487
rect -108 -507 -104 -487
rect 53 -500 57 -460
rect 61 -500 65 -460
rect 83 -500 87 -460
rect 91 -500 95 -460
rect -146 -542 -142 -522
rect -138 -542 -134 -522
rect -116 -542 -112 -522
rect -108 -542 -104 -522
rect 53 -555 57 -515
rect 61 -555 65 -515
rect 83 -555 87 -515
rect 91 -555 95 -515
rect 113 -554 117 -514
rect 121 -554 125 -514
rect 173 -526 177 -506
rect 181 -526 185 -506
rect 610 -339 614 -319
rect 618 -339 622 -319
rect 640 -339 644 -319
rect 648 -339 652 -319
rect 670 -332 674 -312
rect 678 -332 682 -312
rect 610 -374 614 -354
rect 618 -374 622 -354
rect 640 -374 644 -354
rect 648 -374 652 -354
rect 550 -408 554 -388
rect 558 -408 562 -388
rect 580 -408 584 -388
rect 588 -408 592 -388
rect 460 -500 464 -460
rect 468 -500 472 -460
rect 490 -500 494 -460
rect 498 -500 502 -460
rect 520 -500 524 -480
rect 528 -500 532 -480
rect -206 -576 -202 -556
rect -198 -576 -194 -556
rect -176 -576 -172 -556
rect -168 -576 -164 -556
rect 209 -555 213 -515
rect 217 -555 221 -515
rect 269 -527 273 -507
rect 277 -527 281 -507
rect -231 -670 -227 -650
rect -223 -670 -219 -650
rect -141 -677 -137 -657
rect -133 -677 -129 -657
rect -111 -677 -107 -657
rect -103 -677 -99 -657
rect 113 -605 117 -565
rect 121 -605 125 -565
rect 209 -606 213 -566
rect 217 -606 221 -566
rect 460 -555 464 -515
rect 468 -555 472 -515
rect 490 -555 494 -515
rect 498 -555 502 -515
rect 611 -508 615 -488
rect 619 -508 623 -488
rect 641 -508 645 -488
rect 649 -508 653 -488
rect 671 -501 675 -481
rect 679 -501 683 -481
rect 611 -543 615 -523
rect 619 -543 623 -523
rect 641 -543 645 -523
rect 649 -543 653 -523
rect 551 -577 555 -557
rect 559 -577 563 -557
rect 581 -577 585 -557
rect 589 -577 593 -557
rect 317 -657 321 -637
rect 325 -657 329 -637
rect 335 -657 339 -637
rect 343 -657 347 -637
rect 351 -649 355 -629
rect 359 -649 363 -629
rect 521 -671 525 -651
rect 529 -671 533 -651
rect -141 -712 -137 -692
rect -133 -712 -129 -692
rect -111 -712 -107 -692
rect -103 -712 -99 -692
rect -201 -746 -197 -726
rect -193 -746 -189 -726
rect -171 -746 -167 -726
rect -163 -746 -159 -726
rect 616 -678 620 -658
rect 624 -678 628 -658
rect 646 -678 650 -658
rect 654 -678 658 -658
rect 676 -671 680 -651
rect 684 -671 688 -651
rect 616 -713 620 -693
rect 624 -713 628 -693
rect 646 -713 650 -693
rect 654 -713 658 -693
rect 556 -747 560 -727
rect 564 -747 568 -727
rect 586 -747 590 -727
rect 594 -747 598 -727
rect -228 -841 -224 -821
rect -220 -841 -216 -821
rect -138 -848 -134 -828
rect -130 -848 -126 -828
rect -108 -848 -104 -828
rect -100 -848 -96 -828
rect 58 -832 62 -792
rect 66 -832 70 -792
rect 88 -832 92 -792
rect 96 -832 100 -792
rect -138 -883 -134 -863
rect -130 -883 -126 -863
rect -108 -883 -104 -863
rect -100 -883 -96 -863
rect 58 -887 62 -847
rect 66 -887 70 -847
rect 88 -887 92 -847
rect 96 -887 100 -847
rect 461 -831 465 -791
rect 469 -831 473 -791
rect 491 -831 495 -791
rect 499 -831 503 -791
rect -198 -917 -194 -897
rect -190 -917 -186 -897
rect -168 -917 -164 -897
rect -160 -917 -156 -897
rect 317 -910 321 -890
rect 325 -910 329 -890
rect 335 -910 339 -890
rect 343 -910 347 -890
rect 351 -902 355 -882
rect 359 -902 363 -882
rect 461 -886 465 -846
rect 469 -886 473 -846
rect 491 -886 495 -846
rect 499 -886 503 -846
rect -226 -1012 -222 -992
rect -218 -1012 -214 -992
rect -136 -1019 -132 -999
rect -128 -1019 -124 -999
rect -106 -1019 -102 -999
rect -98 -1019 -94 -999
rect -136 -1054 -132 -1034
rect -128 -1054 -124 -1034
rect -106 -1054 -102 -1034
rect -98 -1054 -94 -1034
rect -196 -1088 -192 -1068
rect -188 -1088 -184 -1068
rect -166 -1088 -162 -1068
rect -158 -1088 -154 -1068
rect -223 -1184 -219 -1164
rect -215 -1184 -211 -1164
rect 62 -1165 66 -1125
rect 70 -1165 74 -1125
rect 92 -1165 96 -1125
rect 100 -1165 104 -1125
rect 460 -1162 464 -1122
rect 468 -1162 472 -1122
rect 490 -1162 494 -1122
rect 498 -1162 502 -1122
rect -133 -1191 -129 -1171
rect -125 -1191 -121 -1171
rect -103 -1191 -99 -1171
rect -95 -1191 -91 -1171
rect -133 -1226 -129 -1206
rect -125 -1226 -121 -1206
rect -103 -1226 -99 -1206
rect -95 -1226 -91 -1206
rect 62 -1220 66 -1180
rect 70 -1220 74 -1180
rect 92 -1220 96 -1180
rect 100 -1220 104 -1180
rect 460 -1217 464 -1177
rect 468 -1217 472 -1177
rect 490 -1217 494 -1177
rect 498 -1217 502 -1177
rect -193 -1260 -189 -1240
rect -185 -1260 -181 -1240
rect -163 -1260 -159 -1240
rect -155 -1260 -151 -1240
<< pdcontact >>
rect -238 45 -234 85
rect -230 45 -226 85
rect -208 43 -204 83
rect -200 43 -196 83
rect -178 43 -174 83
rect -170 43 -166 83
rect -148 43 -144 83
rect -140 43 -136 83
rect -118 43 -114 83
rect -110 43 -106 83
rect -88 44 -84 84
rect -80 44 -76 84
rect -54 44 -50 84
rect -46 44 -42 84
rect -23 43 -19 83
rect -15 43 -11 83
rect 11 43 15 83
rect 19 43 23 83
rect -208 -18 -204 22
rect -200 -18 -196 22
rect -178 -18 -174 22
rect -170 -18 -166 22
rect 49 3 53 83
rect 57 3 61 83
rect 79 3 83 83
rect 87 3 91 83
rect 109 43 113 83
rect 117 43 121 83
rect 139 43 143 83
rect 147 43 151 83
rect 169 43 173 83
rect 177 43 181 83
rect 211 43 215 83
rect 219 43 223 83
rect 241 43 245 83
rect 249 43 253 83
rect 271 43 275 83
rect 279 43 283 83
rect -83 -53 -79 -13
rect -75 -53 -71 -13
rect -49 -53 -45 -13
rect -41 -53 -37 -13
rect -18 -54 -14 -14
rect -10 -54 -6 -14
rect 16 -54 20 -14
rect 24 -54 28 -14
rect 317 3 321 83
rect 325 3 329 83
rect 376 43 380 83
rect 384 43 388 83
rect 410 43 414 83
rect 418 43 422 83
rect 459 3 463 83
rect 467 3 471 83
rect 489 3 493 83
rect 497 3 501 83
rect 519 43 523 83
rect 527 43 531 83
rect 549 42 553 82
rect 557 42 561 82
rect 579 42 583 82
rect 587 42 591 82
rect 609 42 613 82
rect 617 42 621 82
rect 639 42 643 82
rect 647 42 651 82
rect 669 43 673 83
rect 677 43 681 83
rect -235 -127 -231 -87
rect -227 -127 -223 -87
rect -205 -128 -201 -88
rect -197 -128 -193 -88
rect -175 -128 -171 -88
rect -167 -128 -163 -88
rect -145 -128 -141 -88
rect -137 -128 -133 -88
rect -115 -128 -111 -88
rect -107 -128 -103 -88
rect 49 -102 53 -22
rect 57 -102 61 -22
rect 79 -102 83 -22
rect 87 -102 91 -22
rect -82 -149 -78 -109
rect -74 -149 -70 -109
rect -48 -149 -44 -109
rect -40 -149 -36 -109
rect -205 -189 -201 -149
rect -197 -189 -193 -149
rect -175 -189 -171 -149
rect -167 -189 -163 -149
rect -17 -150 -13 -110
rect -9 -150 -5 -110
rect 17 -150 21 -110
rect 25 -150 29 -110
rect 109 -135 113 -95
rect 117 -135 121 -95
rect 139 -135 143 -95
rect 147 -135 151 -95
rect 169 -135 173 -95
rect 177 -135 181 -95
rect 212 -135 216 -95
rect 220 -135 224 -95
rect 242 -135 246 -95
rect 250 -135 254 -95
rect 272 -135 276 -95
rect 280 -135 284 -95
rect 317 -108 321 -28
rect 325 -108 329 -28
rect 381 -54 385 -14
rect 389 -54 393 -14
rect 415 -54 419 -14
rect 423 -54 427 -14
rect 549 -19 553 21
rect 557 -19 561 21
rect 579 -19 583 21
rect 587 -19 591 21
rect 351 -107 355 -67
rect 359 -107 363 -67
rect 459 -102 463 -22
rect 467 -102 471 -22
rect 489 -102 493 -22
rect 497 -102 501 -22
rect -77 -246 -73 -206
rect -69 -246 -65 -206
rect -43 -246 -39 -206
rect -35 -246 -31 -206
rect -237 -296 -233 -256
rect -229 -296 -225 -256
rect -207 -297 -203 -257
rect -199 -297 -195 -257
rect -177 -297 -173 -257
rect -169 -297 -165 -257
rect -147 -297 -143 -257
rect -139 -297 -135 -257
rect -117 -297 -113 -257
rect -109 -297 -105 -257
rect -12 -247 -8 -207
rect -4 -247 0 -207
rect 22 -247 26 -207
rect 30 -247 34 -207
rect 382 -150 386 -110
rect 390 -150 394 -110
rect 416 -150 420 -110
rect 424 -150 428 -110
rect 519 -128 523 -88
rect 527 -128 531 -88
rect -207 -358 -203 -318
rect -199 -358 -195 -318
rect -177 -358 -173 -318
rect -169 -358 -165 -318
rect 53 -328 57 -248
rect 61 -328 65 -248
rect 83 -328 87 -248
rect 91 -328 95 -248
rect 317 -250 321 -170
rect 325 -250 329 -170
rect 552 -129 556 -89
rect 560 -129 564 -89
rect 582 -129 586 -89
rect 590 -129 594 -89
rect 612 -129 616 -89
rect 620 -129 624 -89
rect 642 -129 646 -89
rect 650 -129 654 -89
rect 672 -128 676 -88
rect 680 -128 684 -88
rect 387 -247 391 -207
rect 395 -247 399 -207
rect 421 -247 425 -207
rect 429 -247 433 -207
rect 552 -190 556 -150
rect 560 -190 564 -150
rect 582 -190 586 -150
rect 590 -190 594 -150
rect 113 -313 117 -273
rect 121 -313 125 -273
rect 143 -313 147 -273
rect 151 -313 155 -273
rect 173 -313 177 -273
rect 181 -313 185 -273
rect 208 -314 212 -274
rect 216 -314 220 -274
rect 238 -314 242 -274
rect 246 -314 250 -274
rect 268 -314 272 -274
rect 276 -314 280 -274
rect -236 -465 -232 -425
rect -228 -465 -224 -425
rect -206 -466 -202 -426
rect -198 -466 -194 -426
rect -176 -466 -172 -426
rect -168 -466 -164 -426
rect -146 -466 -142 -426
rect -138 -466 -134 -426
rect -116 -466 -112 -426
rect -108 -466 -104 -426
rect 53 -433 57 -353
rect 61 -433 65 -353
rect 83 -433 87 -353
rect 91 -433 95 -353
rect 317 -361 321 -281
rect 325 -361 329 -281
rect 351 -361 355 -321
rect 359 -361 363 -321
rect 460 -328 464 -248
rect 468 -328 472 -248
rect 490 -328 494 -248
rect 498 -328 502 -248
rect 520 -297 524 -257
rect 528 -297 532 -257
rect 550 -298 554 -258
rect 558 -298 562 -258
rect 580 -298 584 -258
rect 588 -298 592 -258
rect 610 -298 614 -258
rect 618 -298 622 -258
rect 640 -298 644 -258
rect 648 -298 652 -258
rect 670 -297 674 -257
rect 678 -297 682 -257
rect -206 -527 -202 -487
rect -198 -527 -194 -487
rect -176 -527 -172 -487
rect -168 -527 -164 -487
rect 113 -491 117 -451
rect 121 -491 125 -451
rect 143 -491 147 -451
rect 151 -491 155 -451
rect 173 -491 177 -451
rect 181 -491 185 -451
rect 209 -492 213 -452
rect 217 -492 221 -452
rect 239 -492 243 -452
rect 247 -492 251 -452
rect 269 -492 273 -452
rect 277 -492 281 -452
rect 317 -503 321 -423
rect 325 -503 329 -423
rect 460 -433 464 -353
rect 468 -433 472 -353
rect 490 -433 494 -353
rect 498 -433 502 -353
rect 550 -359 554 -319
rect 558 -359 562 -319
rect 580 -359 584 -319
rect 588 -359 592 -319
rect 520 -465 524 -425
rect 528 -465 532 -425
rect 551 -467 555 -427
rect 559 -467 563 -427
rect 581 -467 585 -427
rect 589 -467 593 -427
rect 611 -467 615 -427
rect 619 -467 623 -427
rect 641 -467 645 -427
rect 649 -467 653 -427
rect 671 -466 675 -426
rect 679 -466 683 -426
rect -231 -635 -227 -595
rect -223 -635 -219 -595
rect -201 -636 -197 -596
rect -193 -636 -189 -596
rect -171 -636 -167 -596
rect -163 -636 -159 -596
rect -141 -636 -137 -596
rect -133 -636 -129 -596
rect -111 -636 -107 -596
rect -103 -636 -99 -596
rect -201 -697 -197 -657
rect -193 -697 -189 -657
rect -171 -697 -167 -657
rect -163 -697 -159 -657
rect 58 -660 62 -580
rect 66 -660 70 -580
rect 88 -660 92 -580
rect 96 -660 100 -580
rect 317 -614 321 -534
rect 325 -614 329 -534
rect 551 -528 555 -488
rect 559 -528 563 -488
rect 581 -528 585 -488
rect 589 -528 593 -488
rect 351 -614 355 -574
rect 359 -614 363 -574
rect 461 -659 465 -579
rect 469 -659 473 -579
rect 491 -659 495 -579
rect 499 -659 503 -579
rect 521 -636 525 -596
rect 529 -636 533 -596
rect 556 -637 560 -597
rect 564 -637 568 -597
rect 586 -637 590 -597
rect 594 -637 598 -597
rect 616 -637 620 -597
rect 624 -637 628 -597
rect 646 -637 650 -597
rect 654 -637 658 -597
rect 676 -636 680 -596
rect 684 -636 688 -596
rect -228 -806 -224 -766
rect -220 -806 -216 -766
rect 58 -765 62 -685
rect 66 -765 70 -685
rect 88 -765 92 -685
rect 96 -765 100 -685
rect 317 -756 321 -676
rect 325 -756 329 -676
rect -198 -807 -194 -767
rect -190 -807 -186 -767
rect -168 -807 -164 -767
rect -160 -807 -156 -767
rect -138 -807 -134 -767
rect -130 -807 -126 -767
rect -108 -807 -104 -767
rect -100 -807 -96 -767
rect 461 -764 465 -684
rect 469 -764 473 -684
rect 491 -764 495 -684
rect 499 -764 503 -684
rect 556 -698 560 -658
rect 564 -698 568 -658
rect 586 -698 590 -658
rect 594 -698 598 -658
rect -198 -868 -194 -828
rect -190 -868 -186 -828
rect -168 -868 -164 -828
rect -160 -868 -156 -828
rect 317 -867 321 -787
rect 325 -867 329 -787
rect 351 -867 355 -827
rect 359 -867 363 -827
rect -226 -977 -222 -937
rect -218 -977 -214 -937
rect -196 -978 -192 -938
rect -188 -978 -184 -938
rect -166 -978 -162 -938
rect -158 -978 -154 -938
rect -136 -978 -132 -938
rect -128 -978 -124 -938
rect -106 -978 -102 -938
rect -98 -978 -94 -938
rect 62 -993 66 -913
rect 70 -993 74 -913
rect 92 -993 96 -913
rect 100 -993 104 -913
rect 460 -990 464 -910
rect 468 -990 472 -910
rect 490 -990 494 -910
rect 498 -990 502 -910
rect -196 -1039 -192 -999
rect -188 -1039 -184 -999
rect -166 -1039 -162 -999
rect -158 -1039 -154 -999
rect 62 -1098 66 -1018
rect 70 -1098 74 -1018
rect 92 -1098 96 -1018
rect 100 -1098 104 -1018
rect 460 -1095 464 -1015
rect 468 -1095 472 -1015
rect 490 -1095 494 -1015
rect 498 -1095 502 -1015
rect -223 -1149 -219 -1109
rect -215 -1149 -211 -1109
rect -193 -1150 -189 -1110
rect -185 -1150 -181 -1110
rect -163 -1150 -159 -1110
rect -155 -1150 -151 -1110
rect -133 -1150 -129 -1110
rect -125 -1150 -121 -1110
rect -103 -1150 -99 -1110
rect -95 -1150 -91 -1110
rect -193 -1211 -189 -1171
rect -185 -1211 -181 -1171
rect -163 -1211 -159 -1171
rect -155 -1211 -151 -1171
<< polysilicon >>
rect -233 85 -231 88
rect -203 83 -201 86
rect -173 83 -171 86
rect -143 83 -141 86
rect -113 83 -111 86
rect -83 84 -81 87
rect -49 84 -47 87
rect -233 30 -231 45
rect -18 83 -16 86
rect 16 83 18 86
rect 54 83 56 86
rect 84 83 86 86
rect 114 83 116 86
rect 144 83 146 86
rect 174 83 176 86
rect 216 83 218 86
rect 246 83 248 86
rect 276 83 278 86
rect 322 83 324 86
rect 381 83 383 86
rect 415 83 417 86
rect 464 83 466 86
rect 494 83 496 86
rect 524 83 526 86
rect -203 29 -201 43
rect -173 29 -171 43
rect -143 29 -141 43
rect -113 29 -111 43
rect -83 29 -81 44
rect -49 29 -47 44
rect -203 22 -201 25
rect -173 22 -171 25
rect -143 22 -141 25
rect -113 22 -111 25
rect -233 7 -231 10
rect -18 28 -16 43
rect 16 28 18 43
rect -83 6 -81 9
rect -49 6 -47 9
rect -18 5 -16 8
rect 16 5 18 8
rect 114 32 116 43
rect 144 32 146 43
rect 174 28 176 43
rect 216 32 218 43
rect 246 32 248 43
rect 276 28 278 43
rect 114 20 116 27
rect -143 -6 -141 2
rect -113 -6 -111 2
rect 54 -8 56 3
rect 84 -8 86 3
rect -143 -13 -141 -10
rect -113 -13 -111 -10
rect -78 -13 -76 -10
rect -44 -13 -42 -10
rect -203 -29 -201 -18
rect -173 -29 -171 -18
rect -203 -47 -201 -40
rect -173 -47 -171 -40
rect -143 -41 -141 -33
rect -113 -41 -111 -33
rect -13 -14 -11 -11
rect 21 -14 23 -11
rect -203 -70 -201 -67
rect -173 -70 -171 -67
rect -78 -68 -76 -53
rect -44 -68 -42 -53
rect 54 -22 56 -19
rect 84 -22 86 -19
rect 216 20 218 27
rect 174 5 176 8
rect 276 5 278 8
rect 381 28 383 43
rect 415 28 417 43
rect 381 5 383 8
rect 415 5 417 8
rect 554 82 556 85
rect 584 82 586 85
rect 614 82 616 85
rect 644 82 646 85
rect 674 83 676 86
rect 524 28 526 43
rect 554 28 556 42
rect 584 28 586 42
rect 614 28 616 42
rect 644 28 646 42
rect 674 28 676 43
rect 554 21 556 24
rect 584 21 586 24
rect 614 21 616 24
rect 644 21 646 24
rect 524 5 526 8
rect 322 -10 324 3
rect 464 -8 466 3
rect 494 -8 496 3
rect 386 -14 388 -11
rect 420 -14 422 -11
rect -230 -87 -228 -84
rect -200 -88 -198 -85
rect -170 -88 -168 -85
rect -140 -88 -138 -85
rect -110 -88 -108 -85
rect -13 -69 -11 -54
rect 21 -69 23 -54
rect -230 -142 -228 -127
rect -78 -91 -76 -88
rect -44 -91 -42 -88
rect -13 -92 -11 -89
rect 21 -92 23 -89
rect 114 -23 116 -20
rect 216 -23 218 -20
rect 322 -28 324 -15
rect 114 -31 116 -28
rect 216 -31 218 -28
rect 114 -78 116 -71
rect 216 -78 218 -71
rect 114 -95 116 -92
rect 144 -95 146 -92
rect 174 -95 176 -92
rect 217 -95 219 -92
rect 247 -95 249 -92
rect 277 -95 279 -92
rect -77 -109 -75 -106
rect -43 -109 -41 -106
rect -200 -142 -198 -128
rect -170 -142 -168 -128
rect -140 -142 -138 -128
rect -110 -142 -108 -128
rect -200 -149 -198 -146
rect -170 -149 -168 -146
rect -140 -149 -138 -146
rect -110 -149 -108 -146
rect -12 -110 -10 -107
rect 22 -110 24 -107
rect -230 -165 -228 -162
rect -77 -164 -75 -149
rect -43 -164 -41 -149
rect 54 -113 56 -102
rect 84 -113 86 -102
rect 54 -129 56 -122
rect 84 -129 86 -122
rect -140 -177 -138 -169
rect -110 -177 -108 -169
rect -140 -184 -138 -181
rect -110 -184 -108 -181
rect -12 -165 -10 -150
rect 22 -165 24 -150
rect -200 -200 -198 -189
rect -170 -200 -168 -189
rect -77 -187 -75 -184
rect -43 -187 -41 -184
rect 674 5 676 8
rect 614 -7 616 1
rect 644 -7 646 1
rect 614 -14 616 -11
rect 644 -14 646 -11
rect 464 -22 466 -19
rect 494 -22 496 -19
rect 356 -67 358 -64
rect 386 -69 388 -54
rect 420 -69 422 -54
rect 386 -92 388 -89
rect 420 -92 422 -89
rect 554 -30 556 -19
rect 584 -30 586 -19
rect 554 -48 556 -41
rect 584 -48 586 -41
rect 614 -42 616 -34
rect 644 -42 646 -34
rect 554 -71 556 -68
rect 584 -71 586 -68
rect 524 -88 526 -85
rect 322 -118 324 -108
rect 356 -122 358 -107
rect 387 -110 389 -107
rect 421 -110 423 -107
rect 322 -131 324 -124
rect 340 -131 342 -124
rect 114 -146 116 -135
rect 144 -146 146 -135
rect 174 -150 176 -135
rect 217 -146 219 -135
rect 247 -146 249 -135
rect 277 -150 279 -135
rect 114 -158 116 -151
rect 54 -175 56 -169
rect 84 -175 86 -169
rect 54 -184 56 -181
rect 84 -184 86 -181
rect -12 -188 -10 -185
rect 22 -188 24 -185
rect -200 -218 -198 -211
rect -170 -218 -168 -211
rect -140 -212 -138 -204
rect -110 -212 -108 -204
rect -72 -206 -70 -203
rect -38 -206 -36 -203
rect -200 -241 -198 -238
rect -170 -241 -168 -238
rect -7 -207 -5 -204
rect 27 -207 29 -204
rect -232 -256 -230 -253
rect -202 -257 -200 -254
rect -172 -257 -170 -254
rect -142 -257 -140 -254
rect -112 -257 -110 -254
rect -232 -311 -230 -296
rect -72 -261 -70 -246
rect -38 -261 -36 -246
rect 217 -158 219 -151
rect 174 -173 176 -170
rect 356 -145 358 -142
rect 464 -113 466 -102
rect 494 -113 496 -102
rect 464 -129 466 -122
rect 494 -129 496 -122
rect 557 -89 559 -86
rect 587 -89 589 -86
rect 617 -89 619 -86
rect 647 -89 649 -86
rect 677 -88 679 -85
rect 322 -154 324 -151
rect 340 -154 342 -151
rect 387 -165 389 -150
rect 421 -165 423 -150
rect 322 -170 324 -167
rect 277 -173 279 -170
rect 114 -201 116 -198
rect 217 -201 219 -198
rect 114 -209 116 -206
rect 217 -209 219 -206
rect 54 -231 56 -224
rect 84 -231 86 -224
rect -7 -262 -5 -247
rect 27 -262 29 -247
rect 58 -248 60 -245
rect 88 -248 90 -245
rect -72 -284 -70 -281
rect -38 -284 -36 -281
rect -7 -285 -5 -282
rect 27 -285 29 -282
rect -202 -311 -200 -297
rect -172 -311 -170 -297
rect -142 -311 -140 -297
rect -112 -311 -110 -297
rect -202 -318 -200 -315
rect -172 -318 -170 -315
rect -142 -318 -140 -315
rect -112 -318 -110 -315
rect -232 -334 -230 -331
rect 114 -256 116 -249
rect 217 -256 219 -249
rect 524 -143 526 -128
rect 557 -143 559 -129
rect 587 -143 589 -129
rect 617 -143 619 -129
rect 647 -143 649 -129
rect 677 -143 679 -128
rect 557 -150 559 -147
rect 587 -150 589 -147
rect 617 -150 619 -147
rect 647 -150 649 -147
rect 524 -166 526 -163
rect 464 -175 466 -169
rect 494 -175 496 -169
rect 464 -184 466 -181
rect 494 -184 496 -181
rect 387 -188 389 -185
rect 421 -188 423 -185
rect 392 -207 394 -204
rect 426 -207 428 -204
rect 677 -166 679 -163
rect 617 -178 619 -170
rect 647 -178 649 -170
rect 617 -185 619 -182
rect 647 -185 649 -182
rect 557 -201 559 -190
rect 587 -201 589 -190
rect 557 -219 559 -212
rect 587 -219 589 -212
rect 617 -213 619 -205
rect 647 -213 649 -205
rect 464 -231 466 -224
rect 494 -231 496 -224
rect 557 -242 559 -239
rect 587 -242 589 -239
rect 322 -263 324 -250
rect 392 -262 394 -247
rect 426 -262 428 -247
rect 465 -248 467 -245
rect 495 -248 497 -245
rect 118 -273 120 -270
rect 148 -273 150 -270
rect 178 -273 180 -270
rect 213 -274 215 -271
rect 243 -274 245 -271
rect 273 -274 275 -271
rect 118 -324 120 -313
rect 148 -324 150 -313
rect 178 -328 180 -313
rect 322 -281 324 -268
rect 213 -325 215 -314
rect 243 -325 245 -314
rect -142 -346 -140 -338
rect -112 -346 -110 -338
rect 58 -339 60 -328
rect 88 -339 90 -328
rect 118 -336 120 -329
rect -142 -353 -140 -350
rect -112 -353 -110 -350
rect 58 -353 60 -350
rect 88 -353 90 -350
rect -202 -369 -200 -358
rect -172 -369 -170 -358
rect -202 -387 -200 -380
rect -172 -387 -170 -380
rect -142 -381 -140 -373
rect -112 -381 -110 -373
rect -202 -410 -200 -407
rect -172 -410 -170 -407
rect -231 -425 -229 -422
rect -201 -426 -199 -423
rect -171 -426 -169 -423
rect -141 -426 -139 -423
rect -111 -426 -109 -423
rect -231 -480 -229 -465
rect 273 -329 275 -314
rect 213 -337 215 -330
rect 178 -351 180 -348
rect 118 -379 120 -376
rect 273 -352 275 -349
rect 392 -285 394 -282
rect 426 -285 428 -282
rect 356 -321 358 -318
rect 525 -257 527 -254
rect 555 -258 557 -255
rect 585 -258 587 -255
rect 615 -258 617 -255
rect 645 -258 647 -255
rect 675 -257 677 -254
rect 525 -312 527 -297
rect 555 -312 557 -298
rect 585 -312 587 -298
rect 615 -312 617 -298
rect 645 -312 647 -298
rect 675 -312 677 -297
rect 465 -339 467 -328
rect 495 -339 497 -328
rect 555 -319 557 -316
rect 585 -319 587 -316
rect 615 -319 617 -316
rect 645 -319 647 -316
rect 525 -335 527 -332
rect 465 -353 467 -350
rect 495 -353 497 -350
rect 322 -371 324 -361
rect 356 -376 358 -361
rect 213 -380 215 -377
rect 322 -384 324 -377
rect 340 -384 342 -377
rect 118 -387 120 -384
rect 213 -388 215 -385
rect 58 -444 60 -433
rect 88 -444 90 -433
rect 118 -434 120 -427
rect 356 -399 358 -396
rect 322 -407 324 -404
rect 340 -407 342 -404
rect 322 -423 324 -420
rect 213 -435 215 -428
rect 118 -451 120 -448
rect 148 -451 150 -448
rect 178 -451 180 -448
rect 58 -460 60 -453
rect 88 -460 90 -453
rect -201 -480 -199 -466
rect -171 -480 -169 -466
rect -141 -480 -139 -466
rect -111 -480 -109 -466
rect -201 -487 -199 -484
rect -171 -487 -169 -484
rect -141 -487 -139 -484
rect -111 -487 -109 -484
rect -231 -503 -229 -500
rect 214 -452 216 -449
rect 244 -452 246 -449
rect 274 -452 276 -449
rect 58 -506 60 -500
rect 88 -506 90 -500
rect 118 -502 120 -491
rect 148 -502 150 -491
rect 178 -506 180 -491
rect 214 -503 216 -492
rect 244 -503 246 -492
rect -141 -515 -139 -507
rect -111 -515 -109 -507
rect 58 -515 60 -512
rect 88 -515 90 -512
rect 118 -514 120 -507
rect -141 -522 -139 -519
rect -111 -522 -109 -519
rect -201 -538 -199 -527
rect -171 -538 -169 -527
rect -201 -556 -199 -549
rect -171 -556 -169 -549
rect -141 -550 -139 -542
rect -111 -550 -109 -542
rect 274 -507 276 -492
rect 675 -335 677 -332
rect 615 -347 617 -339
rect 645 -347 647 -339
rect 615 -354 617 -351
rect 645 -354 647 -351
rect 555 -370 557 -359
rect 585 -370 587 -359
rect 555 -388 557 -381
rect 585 -388 587 -381
rect 615 -382 617 -374
rect 645 -382 647 -374
rect 555 -411 557 -408
rect 585 -411 587 -408
rect 525 -425 527 -422
rect 465 -444 467 -433
rect 495 -444 497 -433
rect 465 -460 467 -453
rect 495 -460 497 -453
rect 556 -427 558 -424
rect 586 -427 588 -424
rect 616 -427 618 -424
rect 646 -427 648 -424
rect 676 -426 678 -423
rect 525 -480 527 -465
rect 556 -481 558 -467
rect 586 -481 588 -467
rect 616 -481 618 -467
rect 646 -481 648 -467
rect 676 -481 678 -466
rect 556 -488 558 -485
rect 586 -488 588 -485
rect 616 -488 618 -485
rect 646 -488 648 -485
rect 214 -515 216 -508
rect 178 -529 180 -526
rect 58 -562 60 -555
rect 88 -562 90 -555
rect 118 -557 120 -554
rect 322 -516 324 -503
rect 465 -506 467 -500
rect 495 -506 497 -500
rect 525 -503 527 -500
rect 465 -515 467 -512
rect 495 -515 497 -512
rect 274 -530 276 -527
rect 322 -534 324 -521
rect 214 -558 216 -555
rect 118 -565 120 -562
rect -201 -579 -199 -576
rect -171 -579 -169 -576
rect 63 -580 65 -577
rect 93 -580 95 -577
rect -226 -595 -224 -592
rect -196 -596 -194 -593
rect -166 -596 -164 -593
rect -136 -596 -134 -593
rect -106 -596 -104 -593
rect -226 -650 -224 -635
rect -196 -650 -194 -636
rect -166 -650 -164 -636
rect -136 -650 -134 -636
rect -106 -650 -104 -636
rect -196 -657 -194 -654
rect -166 -657 -164 -654
rect -136 -657 -134 -654
rect -106 -657 -104 -654
rect -226 -673 -224 -670
rect 214 -566 216 -563
rect 118 -612 120 -605
rect 214 -613 216 -606
rect 676 -504 678 -501
rect 616 -516 618 -508
rect 646 -516 648 -508
rect 616 -523 618 -520
rect 646 -523 648 -520
rect 556 -539 558 -528
rect 586 -539 588 -528
rect 465 -562 467 -555
rect 495 -562 497 -555
rect 556 -557 558 -550
rect 586 -557 588 -550
rect 616 -551 618 -543
rect 646 -551 648 -543
rect 356 -574 358 -571
rect 466 -579 468 -576
rect 496 -579 498 -576
rect 322 -624 324 -614
rect 356 -629 358 -614
rect 322 -637 324 -630
rect 340 -637 342 -630
rect 356 -652 358 -649
rect 322 -660 324 -657
rect 340 -660 342 -657
rect 556 -580 558 -577
rect 586 -580 588 -577
rect 526 -596 528 -593
rect 561 -597 563 -594
rect 591 -597 593 -594
rect 621 -597 623 -594
rect 651 -597 653 -594
rect 681 -596 683 -593
rect 526 -651 528 -636
rect 561 -651 563 -637
rect 591 -651 593 -637
rect 621 -651 623 -637
rect 651 -651 653 -637
rect 681 -651 683 -636
rect 63 -671 65 -660
rect 93 -671 95 -660
rect 466 -670 468 -659
rect 496 -670 498 -659
rect 561 -658 563 -655
rect 591 -658 593 -655
rect 621 -658 623 -655
rect 651 -658 653 -655
rect 322 -676 324 -673
rect 526 -674 528 -671
rect -136 -685 -134 -677
rect -106 -685 -104 -677
rect 63 -685 65 -682
rect 93 -685 95 -682
rect -136 -692 -134 -689
rect -106 -692 -104 -689
rect -196 -708 -194 -697
rect -166 -708 -164 -697
rect -196 -726 -194 -719
rect -166 -726 -164 -719
rect -136 -720 -134 -712
rect -106 -720 -104 -712
rect -196 -749 -194 -746
rect -166 -749 -164 -746
rect -223 -766 -221 -763
rect -193 -767 -191 -764
rect -163 -767 -161 -764
rect -133 -767 -131 -764
rect -103 -767 -101 -764
rect 466 -684 468 -681
rect 496 -684 498 -681
rect -223 -821 -221 -806
rect 63 -776 65 -765
rect 93 -776 95 -765
rect 322 -769 324 -756
rect 681 -674 683 -671
rect 621 -686 623 -678
rect 651 -686 653 -678
rect 621 -693 623 -690
rect 651 -693 653 -690
rect 561 -709 563 -698
rect 591 -709 593 -698
rect 561 -727 563 -720
rect 591 -727 593 -720
rect 621 -721 623 -713
rect 651 -721 653 -713
rect 561 -750 563 -747
rect 591 -750 593 -747
rect 63 -792 65 -785
rect 93 -792 95 -785
rect 322 -787 324 -774
rect 466 -775 468 -764
rect 496 -775 498 -764
rect -193 -821 -191 -807
rect -163 -821 -161 -807
rect -133 -821 -131 -807
rect -103 -821 -101 -807
rect -193 -828 -191 -825
rect -163 -828 -161 -825
rect -133 -828 -131 -825
rect -103 -828 -101 -825
rect -223 -844 -221 -841
rect 63 -838 65 -832
rect 93 -838 95 -832
rect 63 -847 65 -844
rect 93 -847 95 -844
rect -133 -856 -131 -848
rect -103 -856 -101 -848
rect -133 -863 -131 -860
rect -103 -863 -101 -860
rect -193 -879 -191 -868
rect -163 -879 -161 -868
rect -193 -897 -191 -890
rect -163 -897 -161 -890
rect -133 -891 -131 -883
rect -103 -891 -101 -883
rect 466 -791 468 -784
rect 496 -791 498 -784
rect 356 -827 358 -824
rect 466 -837 468 -831
rect 496 -837 498 -831
rect 466 -846 468 -843
rect 496 -846 498 -843
rect 322 -877 324 -867
rect 356 -882 358 -867
rect 63 -894 65 -887
rect 93 -894 95 -887
rect 322 -890 324 -883
rect 340 -890 342 -883
rect 466 -893 468 -886
rect 496 -893 498 -886
rect 356 -905 358 -902
rect 465 -910 467 -907
rect 495 -910 497 -907
rect 67 -913 69 -910
rect 97 -913 99 -910
rect 322 -913 324 -910
rect 340 -913 342 -910
rect -193 -920 -191 -917
rect -163 -920 -161 -917
rect -221 -937 -219 -934
rect -191 -938 -189 -935
rect -161 -938 -159 -935
rect -131 -938 -129 -935
rect -101 -938 -99 -935
rect -221 -992 -219 -977
rect -191 -992 -189 -978
rect -161 -992 -159 -978
rect -131 -992 -129 -978
rect -101 -992 -99 -978
rect -191 -999 -189 -996
rect -161 -999 -159 -996
rect -131 -999 -129 -996
rect -101 -999 -99 -996
rect -221 -1015 -219 -1012
rect 67 -1004 69 -993
rect 97 -1004 99 -993
rect 465 -1001 467 -990
rect 495 -1001 497 -990
rect 465 -1015 467 -1012
rect 495 -1015 497 -1012
rect 67 -1018 69 -1015
rect 97 -1018 99 -1015
rect -131 -1027 -129 -1019
rect -101 -1027 -99 -1019
rect -131 -1034 -129 -1031
rect -101 -1034 -99 -1031
rect -191 -1050 -189 -1039
rect -161 -1050 -159 -1039
rect -191 -1068 -189 -1061
rect -161 -1068 -159 -1061
rect -131 -1062 -129 -1054
rect -101 -1062 -99 -1054
rect -191 -1091 -189 -1088
rect -161 -1091 -159 -1088
rect -218 -1109 -216 -1106
rect -188 -1110 -186 -1107
rect -158 -1110 -156 -1107
rect -128 -1110 -126 -1107
rect -98 -1110 -96 -1107
rect 67 -1109 69 -1098
rect 97 -1109 99 -1098
rect 465 -1106 467 -1095
rect 495 -1106 497 -1095
rect -218 -1164 -216 -1149
rect 67 -1125 69 -1118
rect 97 -1125 99 -1118
rect 465 -1122 467 -1115
rect 495 -1122 497 -1115
rect -188 -1164 -186 -1150
rect -158 -1164 -156 -1150
rect -128 -1164 -126 -1150
rect -98 -1164 -96 -1150
rect -188 -1171 -186 -1168
rect -158 -1171 -156 -1168
rect -128 -1171 -126 -1168
rect -98 -1171 -96 -1168
rect 67 -1171 69 -1165
rect 97 -1171 99 -1165
rect 465 -1168 467 -1162
rect 495 -1168 497 -1162
rect -218 -1187 -216 -1184
rect 465 -1177 467 -1174
rect 495 -1177 497 -1174
rect 67 -1180 69 -1177
rect 97 -1180 99 -1177
rect -128 -1199 -126 -1191
rect -98 -1199 -96 -1191
rect -128 -1206 -126 -1203
rect -98 -1206 -96 -1203
rect -188 -1222 -186 -1211
rect -158 -1222 -156 -1211
rect -188 -1240 -186 -1233
rect -158 -1240 -156 -1233
rect -128 -1234 -126 -1226
rect -98 -1234 -96 -1226
rect 67 -1227 69 -1220
rect 97 -1227 99 -1220
rect 465 -1224 467 -1217
rect 495 -1224 497 -1217
rect -188 -1263 -186 -1260
rect -158 -1263 -156 -1260
<< polycontact >>
rect -237 33 -233 37
rect -207 29 -203 33
rect -177 29 -173 33
rect -147 29 -143 33
rect -117 29 -113 33
rect -87 32 -83 36
rect -53 32 -49 36
rect -22 31 -18 35
rect 12 31 16 35
rect 110 32 114 36
rect 140 32 144 36
rect 170 31 174 35
rect 212 32 216 36
rect 242 32 246 36
rect 272 31 276 35
rect 110 23 114 27
rect -141 -6 -137 -2
rect -111 -6 -107 -2
rect 50 -8 54 -4
rect 80 -8 84 -4
rect -201 -29 -197 -25
rect -171 -29 -167 -25
rect -201 -44 -197 -40
rect -171 -44 -167 -40
rect -147 -41 -143 -37
rect -117 -41 -113 -37
rect -82 -65 -78 -61
rect -48 -65 -44 -61
rect 212 23 216 27
rect 377 31 381 35
rect 411 31 415 35
rect 520 31 524 35
rect 550 28 554 32
rect 580 28 584 32
rect 610 28 614 32
rect 640 28 644 32
rect 670 31 674 35
rect 324 -10 328 -6
rect 460 -8 464 -4
rect 490 -8 494 -4
rect -17 -66 -13 -62
rect 17 -66 21 -62
rect -234 -139 -230 -135
rect 324 -19 328 -15
rect 110 -78 114 -74
rect 212 -78 216 -74
rect -204 -142 -200 -138
rect -174 -142 -170 -138
rect -144 -142 -140 -138
rect -114 -142 -110 -138
rect -81 -161 -77 -157
rect -47 -161 -43 -157
rect 56 -113 60 -109
rect 86 -113 90 -109
rect 56 -126 60 -122
rect 86 -126 90 -122
rect -16 -162 -12 -158
rect -138 -177 -134 -173
rect -108 -177 -104 -173
rect 18 -162 22 -158
rect -198 -200 -194 -196
rect -168 -200 -164 -196
rect 616 -7 620 -3
rect 646 -7 650 -3
rect 382 -66 386 -62
rect 416 -66 420 -62
rect 556 -30 560 -26
rect 586 -30 590 -26
rect 556 -45 560 -41
rect 586 -45 590 -41
rect 610 -42 614 -38
rect 640 -42 644 -38
rect 352 -119 356 -115
rect 318 -128 322 -124
rect 342 -128 346 -124
rect 110 -146 114 -142
rect 140 -146 144 -142
rect 170 -147 174 -143
rect 213 -146 217 -142
rect 243 -146 247 -142
rect 273 -147 277 -143
rect 110 -155 114 -151
rect -198 -215 -194 -211
rect -168 -215 -164 -211
rect -144 -212 -140 -208
rect -114 -212 -110 -208
rect -236 -308 -232 -304
rect -76 -258 -72 -254
rect -42 -258 -38 -254
rect 213 -155 217 -151
rect 466 -113 470 -109
rect 496 -113 500 -109
rect 466 -126 470 -122
rect 496 -126 500 -122
rect 383 -162 387 -158
rect 417 -162 421 -158
rect 56 -231 60 -227
rect 86 -231 90 -227
rect -11 -259 -7 -255
rect 23 -259 27 -255
rect -206 -311 -202 -307
rect -176 -311 -172 -307
rect -146 -311 -142 -307
rect -116 -311 -112 -307
rect 110 -256 114 -252
rect 213 -256 217 -252
rect 520 -140 524 -136
rect 553 -143 557 -139
rect 583 -143 587 -139
rect 613 -143 617 -139
rect 643 -143 647 -139
rect 673 -140 677 -136
rect 619 -178 623 -174
rect 649 -178 653 -174
rect 559 -201 563 -197
rect 589 -201 593 -197
rect 559 -216 563 -212
rect 589 -216 593 -212
rect 613 -213 617 -209
rect 643 -213 647 -209
rect 466 -231 470 -227
rect 496 -231 500 -227
rect 388 -259 392 -255
rect 324 -263 328 -259
rect 422 -259 426 -255
rect 114 -324 118 -320
rect 144 -324 148 -320
rect 174 -325 178 -321
rect 324 -272 328 -268
rect 209 -325 213 -321
rect 239 -325 243 -321
rect 269 -326 273 -322
rect -140 -346 -136 -342
rect 54 -339 58 -335
rect 84 -339 88 -335
rect 114 -333 118 -329
rect -110 -346 -106 -342
rect -200 -369 -196 -365
rect -170 -369 -166 -365
rect -200 -384 -196 -380
rect -170 -384 -166 -380
rect -146 -381 -142 -377
rect -116 -381 -112 -377
rect -235 -477 -231 -473
rect 209 -334 213 -330
rect 521 -309 525 -305
rect 551 -312 555 -308
rect 581 -312 585 -308
rect 611 -312 615 -308
rect 641 -312 645 -308
rect 671 -309 675 -305
rect 461 -339 465 -335
rect 491 -339 495 -335
rect 352 -373 356 -369
rect 318 -381 322 -377
rect 342 -381 346 -377
rect 60 -444 64 -440
rect 114 -434 118 -430
rect 209 -435 213 -431
rect 90 -444 94 -440
rect 60 -457 64 -453
rect 90 -457 94 -453
rect -205 -480 -201 -476
rect -175 -480 -171 -476
rect -145 -480 -141 -476
rect -115 -480 -111 -476
rect 114 -502 118 -498
rect 144 -502 148 -498
rect 174 -503 178 -499
rect 210 -503 214 -499
rect 240 -503 244 -499
rect 270 -504 274 -500
rect -139 -515 -135 -511
rect 114 -511 118 -507
rect -109 -515 -105 -511
rect -199 -538 -195 -534
rect -169 -538 -165 -534
rect -199 -553 -195 -549
rect -169 -553 -165 -549
rect -145 -550 -141 -546
rect -115 -550 -111 -546
rect 617 -347 621 -343
rect 647 -347 651 -343
rect 557 -370 561 -366
rect 587 -370 591 -366
rect 557 -385 561 -381
rect 587 -385 591 -381
rect 611 -382 615 -378
rect 641 -382 645 -378
rect 467 -444 471 -440
rect 497 -444 501 -440
rect 467 -457 471 -453
rect 497 -457 501 -453
rect 521 -477 525 -473
rect 552 -481 556 -477
rect 582 -481 586 -477
rect 612 -481 616 -477
rect 642 -481 646 -477
rect 672 -478 676 -474
rect 210 -512 214 -508
rect 60 -562 64 -558
rect 324 -516 328 -512
rect 324 -525 328 -521
rect 90 -562 94 -558
rect -230 -647 -226 -643
rect -200 -650 -196 -646
rect -170 -650 -166 -646
rect -140 -650 -136 -646
rect -110 -650 -106 -646
rect 114 -612 118 -608
rect 210 -613 214 -609
rect 618 -516 622 -512
rect 648 -516 652 -512
rect 558 -539 562 -535
rect 588 -539 592 -535
rect 467 -562 471 -558
rect 558 -554 562 -550
rect 588 -554 592 -550
rect 612 -551 616 -547
rect 642 -551 646 -547
rect 497 -562 501 -558
rect 352 -626 356 -622
rect 318 -634 322 -630
rect 342 -634 346 -630
rect 522 -648 526 -644
rect 557 -651 561 -647
rect 587 -651 591 -647
rect 617 -651 621 -647
rect 647 -651 651 -647
rect 677 -648 681 -644
rect 59 -671 63 -667
rect 89 -671 93 -667
rect 462 -670 466 -666
rect 492 -670 496 -666
rect -134 -685 -130 -681
rect -104 -685 -100 -681
rect -194 -708 -190 -704
rect -164 -708 -160 -704
rect -194 -723 -190 -719
rect -164 -723 -160 -719
rect -140 -720 -136 -716
rect -110 -720 -106 -716
rect -227 -818 -223 -814
rect 65 -776 69 -772
rect 623 -686 627 -682
rect 653 -686 657 -682
rect 563 -709 567 -705
rect 593 -709 597 -705
rect 563 -724 567 -720
rect 593 -724 597 -720
rect 617 -721 621 -717
rect 647 -721 651 -717
rect 324 -769 328 -765
rect 95 -776 99 -772
rect 65 -789 69 -785
rect 95 -789 99 -785
rect 324 -778 328 -774
rect 468 -775 472 -771
rect 498 -775 502 -771
rect -197 -821 -193 -817
rect -167 -821 -163 -817
rect -137 -821 -133 -817
rect -107 -821 -103 -817
rect -131 -856 -127 -852
rect -101 -856 -97 -852
rect -191 -879 -187 -875
rect -161 -879 -157 -875
rect -191 -894 -187 -890
rect -161 -894 -157 -890
rect -137 -891 -133 -887
rect -107 -891 -103 -887
rect 468 -788 472 -784
rect 498 -788 502 -784
rect 352 -879 356 -875
rect 318 -887 322 -883
rect 65 -894 69 -890
rect 342 -887 346 -883
rect 95 -894 99 -890
rect 468 -893 472 -889
rect 498 -893 502 -889
rect -225 -989 -221 -985
rect -195 -992 -191 -988
rect -165 -992 -161 -988
rect -135 -992 -131 -988
rect -105 -992 -101 -988
rect 63 -1004 67 -1000
rect 93 -1004 97 -1000
rect 461 -1001 465 -997
rect 491 -1001 495 -997
rect -129 -1027 -125 -1023
rect -99 -1027 -95 -1023
rect -189 -1050 -185 -1046
rect -159 -1050 -155 -1046
rect -189 -1065 -185 -1061
rect -159 -1065 -155 -1061
rect -135 -1062 -131 -1058
rect -105 -1062 -101 -1058
rect 69 -1109 73 -1105
rect 99 -1109 103 -1105
rect 467 -1106 471 -1102
rect 497 -1106 501 -1102
rect -222 -1161 -218 -1157
rect 69 -1122 73 -1118
rect 99 -1122 103 -1118
rect 467 -1119 471 -1115
rect 497 -1119 501 -1115
rect -192 -1164 -188 -1160
rect -162 -1164 -158 -1160
rect -132 -1164 -128 -1160
rect -102 -1164 -98 -1160
rect -126 -1199 -122 -1195
rect -96 -1199 -92 -1195
rect -186 -1222 -182 -1218
rect -156 -1222 -152 -1218
rect -186 -1237 -182 -1233
rect -156 -1237 -152 -1233
rect -132 -1234 -128 -1230
rect -102 -1234 -98 -1230
rect 69 -1227 73 -1223
rect 99 -1227 103 -1223
rect 467 -1224 471 -1220
rect 497 -1224 501 -1220
<< metal1 >>
rect -244 89 -220 93
rect -214 89 -190 92
rect -184 89 -160 92
rect -154 89 -130 92
rect -124 89 -100 92
rect -238 85 -234 89
rect -230 37 -226 45
rect -208 83 -204 89
rect -178 83 -174 89
rect -148 83 -144 89
rect -118 83 -114 89
rect -94 88 -70 92
rect -60 88 -36 92
rect -88 84 -84 88
rect -54 84 -50 88
rect -29 87 -5 91
rect 5 87 29 91
rect 43 87 67 91
rect 73 87 97 91
rect 103 87 157 91
rect 163 87 187 91
rect 205 87 259 91
rect 265 87 289 91
rect 311 87 335 91
rect 370 87 394 91
rect 404 87 428 91
rect 453 87 477 91
rect 483 87 507 91
rect 513 87 537 91
rect 543 88 567 91
rect 573 88 597 91
rect 603 88 627 91
rect 633 88 657 91
rect -241 33 -237 37
rect -230 33 -221 37
rect -230 30 -226 33
rect -210 29 -207 33
rect -200 22 -196 43
rect -180 29 -177 33
rect -170 22 -166 43
rect -150 29 -147 33
rect -140 22 -136 43
rect -120 29 -117 33
rect -110 22 -106 43
rect -80 36 -76 44
rect -46 36 -42 44
rect -23 83 -19 87
rect 11 83 15 87
rect 49 83 53 87
rect 79 83 83 87
rect 109 83 113 87
rect 139 83 143 87
rect 169 83 173 87
rect 211 83 215 87
rect 241 83 245 87
rect 271 83 275 87
rect 325 83 329 87
rect -91 32 -87 36
rect -80 32 -71 36
rect -57 32 -53 36
rect -46 32 -38 36
rect -15 35 -11 43
rect 19 35 23 43
rect -80 29 -76 32
rect -46 29 -42 32
rect -26 31 -22 35
rect -15 31 -6 35
rect 8 31 12 35
rect 19 31 27 35
rect -238 5 -234 10
rect -238 1 -226 5
rect -15 28 -11 31
rect 19 28 23 31
rect -88 4 -84 9
rect -54 4 -50 9
rect -148 -13 -144 2
rect -137 -6 -134 -2
rect -118 -13 -114 2
rect -88 0 -76 4
rect -54 0 -42 4
rect -23 3 -19 8
rect 11 3 15 8
rect 108 32 110 36
rect 117 29 121 43
rect 138 32 140 36
rect 147 35 151 43
rect 177 35 181 43
rect 147 31 170 35
rect 177 31 186 35
rect 210 32 212 36
rect 147 29 151 31
rect 108 23 110 27
rect 117 26 151 29
rect 177 28 181 31
rect 117 20 121 26
rect -23 -1 -11 3
rect 11 -1 23 3
rect -107 -6 -104 -2
rect -89 -9 -65 -5
rect -55 -9 -31 -5
rect -83 -13 -79 -9
rect -49 -13 -45 -9
rect -24 -10 0 -6
rect 10 -10 34 -6
rect 48 -8 50 -4
rect -208 -47 -204 -18
rect -197 -29 -193 -25
rect -197 -44 -193 -40
rect -178 -47 -174 -18
rect -167 -29 -163 -25
rect -167 -44 -161 -40
rect -150 -41 -147 -37
rect -140 -44 -136 -33
rect -120 -41 -117 -37
rect -110 -44 -106 -33
rect -150 -47 -136 -44
rect -120 -47 -106 -44
rect -75 -61 -71 -53
rect -41 -61 -37 -53
rect -18 -14 -14 -10
rect 16 -14 20 -10
rect 57 -11 61 3
rect 78 -8 80 -4
rect 87 -11 91 3
rect 57 -14 91 -11
rect 57 -22 61 -14
rect 87 -22 91 -14
rect -86 -65 -82 -61
rect -75 -65 -67 -61
rect -52 -65 -48 -61
rect -41 -65 -33 -61
rect -10 -62 -6 -54
rect 24 -62 28 -54
rect -200 -71 -196 -67
rect -170 -71 -166 -67
rect -75 -68 -71 -65
rect -41 -68 -37 -65
rect -21 -66 -17 -62
rect -10 -66 -2 -62
rect 13 -66 17 -62
rect 24 -66 32 -62
rect -208 -74 -196 -71
rect -178 -74 -166 -71
rect -241 -83 -217 -79
rect -211 -82 -187 -79
rect -181 -82 -157 -79
rect -151 -82 -127 -79
rect -121 -82 -97 -79
rect -235 -87 -231 -83
rect -227 -135 -223 -127
rect -205 -88 -201 -82
rect -175 -88 -171 -82
rect -145 -88 -141 -82
rect -115 -88 -111 -82
rect -10 -69 -6 -66
rect 24 -69 28 -66
rect -83 -93 -79 -88
rect -49 -93 -45 -88
rect -83 -97 -71 -93
rect -49 -97 -37 -93
rect -18 -94 -14 -89
rect 16 -94 20 -89
rect -18 -98 -6 -94
rect 16 -98 28 -94
rect -88 -105 -64 -101
rect -54 -105 -30 -101
rect 219 29 223 43
rect 240 32 242 36
rect 249 35 253 43
rect 279 35 283 43
rect 249 31 272 35
rect 279 31 288 35
rect 249 29 253 31
rect 210 23 212 27
rect 219 26 253 29
rect 279 28 283 31
rect 219 20 223 26
rect 169 3 173 8
rect 169 -1 181 3
rect 271 3 275 8
rect 376 83 380 87
rect 410 83 414 87
rect 459 83 463 87
rect 489 83 493 87
rect 519 83 523 87
rect 384 35 388 43
rect 418 35 422 43
rect 373 31 377 35
rect 384 31 393 35
rect 407 31 411 35
rect 418 31 426 35
rect 384 28 388 31
rect 418 28 422 31
rect 376 3 380 8
rect 410 3 414 8
rect 527 35 531 43
rect 549 82 553 88
rect 579 82 583 88
rect 609 82 613 88
rect 639 82 643 88
rect 663 87 687 91
rect 669 83 673 87
rect 516 31 520 35
rect 527 31 536 35
rect 527 28 531 31
rect 547 28 550 32
rect 271 -1 283 3
rect 109 -31 113 -20
rect 211 -31 215 -20
rect 317 -28 321 3
rect 376 -1 388 3
rect 410 -1 422 3
rect 328 -10 330 -6
rect 375 -10 399 -6
rect 409 -10 433 -6
rect 458 -8 460 -4
rect 381 -14 385 -10
rect 415 -14 419 -10
rect 467 -11 471 3
rect 488 -8 490 -4
rect 497 -11 501 3
rect 557 21 561 42
rect 577 28 580 32
rect 587 21 591 42
rect 607 28 610 32
rect 617 21 621 42
rect 637 28 640 32
rect 647 31 651 42
rect 677 35 681 43
rect 663 31 670 35
rect 677 31 686 35
rect 647 27 666 31
rect 677 28 681 31
rect 647 21 651 27
rect 519 3 523 8
rect 519 -1 531 3
rect 467 -14 501 -11
rect 328 -19 330 -15
rect 108 -78 110 -74
rect 117 -81 121 -71
rect 210 -78 212 -74
rect 219 -81 223 -71
rect 108 -84 121 -81
rect 210 -84 223 -81
rect 103 -91 157 -87
rect 163 -91 187 -87
rect 206 -91 260 -87
rect 266 -91 290 -87
rect 109 -95 113 -91
rect 139 -95 143 -91
rect 169 -95 173 -91
rect 212 -95 216 -91
rect 242 -95 246 -91
rect 272 -95 276 -91
rect -238 -139 -234 -135
rect -227 -139 -218 -135
rect -227 -142 -223 -139
rect -207 -142 -204 -138
rect -197 -149 -193 -128
rect -177 -142 -174 -138
rect -167 -149 -163 -128
rect -147 -142 -144 -138
rect -137 -149 -133 -128
rect -117 -142 -114 -138
rect -107 -149 -103 -128
rect -82 -109 -78 -105
rect -48 -109 -44 -105
rect -23 -106 1 -102
rect 11 -106 35 -102
rect -235 -167 -231 -162
rect -235 -170 -223 -167
rect -74 -157 -70 -149
rect -40 -157 -36 -149
rect -17 -110 -13 -106
rect 17 -110 21 -106
rect -85 -161 -81 -157
rect -74 -161 -65 -157
rect -51 -161 -47 -157
rect -40 -161 -32 -157
rect -9 -158 -5 -150
rect 25 -158 29 -150
rect 49 -116 53 -102
rect 60 -113 62 -109
rect 79 -116 83 -102
rect 90 -113 92 -109
rect 49 -119 83 -116
rect 49 -129 53 -119
rect 60 -126 62 -122
rect 79 -129 83 -119
rect 90 -126 92 -122
rect -74 -164 -70 -161
rect -40 -164 -36 -161
rect -20 -162 -16 -158
rect -9 -162 0 -158
rect 14 -162 18 -158
rect 25 -162 33 -158
rect -145 -184 -141 -169
rect -134 -177 -131 -173
rect -115 -184 -111 -169
rect -104 -177 -101 -173
rect -9 -165 -5 -162
rect 25 -165 29 -162
rect -205 -218 -201 -189
rect -194 -200 -190 -196
rect -194 -215 -190 -211
rect -175 -218 -171 -189
rect -164 -200 -160 -196
rect -82 -189 -78 -184
rect -48 -189 -44 -184
rect 467 -22 471 -14
rect 497 -22 501 -14
rect 345 -63 369 -59
rect 389 -62 393 -54
rect 423 -62 427 -54
rect 351 -67 355 -63
rect 378 -66 382 -62
rect 389 -66 397 -62
rect 412 -66 416 -62
rect 423 -66 431 -62
rect 389 -69 393 -66
rect 423 -69 427 -66
rect 381 -94 385 -89
rect 415 -94 419 -89
rect 381 -98 393 -94
rect 415 -98 427 -94
rect 669 3 673 8
rect 609 -14 613 1
rect 620 -7 623 -3
rect 639 -14 643 1
rect 669 -1 681 3
rect 650 -7 653 -3
rect 549 -48 553 -19
rect 560 -30 564 -26
rect 560 -45 564 -41
rect 579 -48 583 -19
rect 590 -30 594 -26
rect 590 -45 596 -41
rect 607 -42 610 -38
rect 617 -45 621 -34
rect 637 -42 640 -38
rect 647 -45 651 -34
rect 607 -48 621 -45
rect 637 -48 651 -45
rect 557 -72 561 -68
rect 587 -72 591 -68
rect 549 -75 561 -72
rect 579 -75 591 -72
rect 513 -84 537 -80
rect 546 -83 570 -80
rect 576 -83 600 -80
rect 606 -83 630 -80
rect 636 -83 660 -80
rect 519 -88 523 -84
rect 376 -106 400 -102
rect 410 -106 434 -102
rect 325 -115 329 -108
rect 359 -115 363 -107
rect 382 -110 386 -106
rect 416 -110 420 -106
rect 325 -119 352 -115
rect 359 -119 368 -115
rect 325 -124 329 -119
rect 359 -122 363 -119
rect 316 -128 318 -124
rect 325 -127 339 -124
rect 325 -131 329 -127
rect 108 -146 110 -142
rect 117 -149 121 -135
rect 138 -146 140 -142
rect 147 -143 151 -135
rect 177 -143 181 -135
rect 147 -147 170 -143
rect 177 -147 186 -143
rect 211 -146 213 -142
rect 147 -149 151 -147
rect 108 -155 110 -151
rect 117 -152 151 -149
rect 177 -150 181 -147
rect 117 -158 121 -152
rect 57 -184 61 -169
rect 87 -184 91 -169
rect -82 -193 -70 -189
rect -48 -193 -36 -189
rect -17 -190 -13 -185
rect 17 -190 21 -185
rect -17 -194 -5 -190
rect 17 -194 29 -190
rect -83 -202 -59 -198
rect -49 -202 -25 -198
rect -164 -215 -158 -211
rect -147 -212 -144 -208
rect -137 -215 -133 -204
rect -117 -212 -114 -208
rect -107 -215 -103 -204
rect -147 -219 -133 -215
rect -117 -219 -103 -215
rect -77 -206 -73 -202
rect -43 -206 -39 -202
rect -18 -203 6 -199
rect 16 -203 40 -199
rect -197 -242 -193 -238
rect -167 -242 -163 -238
rect -205 -245 -193 -242
rect -175 -245 -163 -242
rect -243 -252 -219 -248
rect -213 -251 -189 -248
rect -183 -251 -159 -248
rect -153 -251 -129 -248
rect -123 -251 -99 -248
rect -237 -256 -233 -252
rect -229 -304 -225 -296
rect -207 -257 -203 -251
rect -177 -257 -173 -251
rect -147 -257 -143 -251
rect -117 -257 -113 -251
rect -69 -254 -65 -246
rect -35 -254 -31 -246
rect -12 -207 -8 -203
rect 22 -207 26 -203
rect 220 -149 224 -135
rect 241 -146 243 -142
rect 250 -143 254 -135
rect 280 -143 284 -135
rect 250 -147 273 -143
rect 280 -147 289 -143
rect 250 -149 254 -147
rect 211 -155 213 -151
rect 220 -152 254 -149
rect 280 -150 284 -147
rect 220 -158 224 -152
rect 169 -175 173 -170
rect 169 -179 181 -175
rect 335 -131 339 -127
rect 346 -128 348 -124
rect 351 -147 355 -142
rect 351 -151 363 -147
rect 317 -155 321 -151
rect 343 -155 347 -151
rect 317 -158 347 -155
rect 390 -158 394 -150
rect 424 -158 428 -150
rect 459 -116 463 -102
rect 470 -113 472 -109
rect 489 -116 493 -102
rect 500 -113 502 -109
rect 459 -119 493 -116
rect 459 -129 463 -119
rect 470 -126 472 -122
rect 489 -129 493 -119
rect 500 -126 502 -122
rect 379 -162 383 -158
rect 390 -162 399 -158
rect 413 -162 417 -158
rect 424 -162 432 -158
rect 311 -166 335 -162
rect 390 -165 394 -162
rect 424 -165 428 -162
rect 325 -170 329 -166
rect 272 -175 276 -170
rect 272 -179 284 -175
rect 109 -209 113 -198
rect 212 -209 216 -198
rect 49 -234 53 -224
rect 60 -231 62 -227
rect 79 -234 83 -224
rect 90 -231 92 -227
rect 49 -237 58 -234
rect 79 -237 88 -234
rect 47 -244 71 -240
rect 77 -244 101 -240
rect -80 -258 -76 -254
rect -69 -258 -61 -254
rect -46 -258 -42 -254
rect -35 -258 -27 -254
rect -4 -255 0 -247
rect 30 -255 34 -247
rect 53 -248 57 -244
rect 83 -248 87 -244
rect -69 -261 -65 -258
rect -35 -261 -31 -258
rect -15 -259 -11 -255
rect -4 -259 4 -255
rect 19 -259 23 -255
rect 30 -259 38 -255
rect -4 -262 0 -259
rect 30 -262 34 -259
rect -77 -286 -73 -281
rect -43 -286 -39 -281
rect -77 -290 -65 -286
rect -43 -290 -31 -286
rect -12 -287 -8 -282
rect 22 -287 26 -282
rect -12 -291 0 -287
rect 22 -291 34 -287
rect -240 -308 -236 -304
rect -229 -308 -220 -304
rect -229 -311 -225 -308
rect -209 -311 -206 -307
rect -199 -318 -195 -297
rect -179 -311 -176 -307
rect -169 -318 -165 -297
rect -149 -311 -146 -307
rect -139 -318 -135 -297
rect -119 -311 -116 -307
rect -109 -318 -105 -297
rect -237 -336 -233 -331
rect -237 -340 -225 -336
rect 108 -256 110 -252
rect 117 -259 121 -249
rect 211 -256 213 -252
rect 220 -259 224 -249
rect 108 -262 121 -259
rect 215 -262 224 -259
rect 527 -136 531 -128
rect 552 -89 556 -83
rect 582 -89 586 -83
rect 612 -89 616 -83
rect 642 -89 646 -83
rect 666 -84 690 -80
rect 672 -88 676 -84
rect 516 -140 520 -136
rect 527 -140 536 -136
rect 527 -143 531 -140
rect 550 -143 553 -139
rect 467 -184 471 -169
rect 497 -184 501 -169
rect 560 -150 564 -129
rect 580 -143 583 -139
rect 590 -150 594 -129
rect 610 -143 613 -139
rect 620 -150 624 -129
rect 640 -143 643 -139
rect 650 -140 654 -129
rect 680 -136 684 -128
rect 666 -140 673 -136
rect 680 -140 689 -136
rect 650 -143 669 -140
rect 680 -143 684 -140
rect 650 -150 654 -143
rect 519 -168 523 -163
rect 519 -172 531 -168
rect 382 -190 386 -185
rect 416 -190 420 -185
rect 382 -194 394 -190
rect 416 -194 428 -190
rect 381 -203 405 -199
rect 415 -203 439 -199
rect 387 -207 391 -203
rect 421 -207 425 -203
rect 672 -168 676 -163
rect 612 -185 616 -170
rect 623 -178 626 -174
rect 642 -185 646 -170
rect 672 -172 684 -168
rect 653 -178 656 -174
rect 552 -219 556 -190
rect 563 -201 567 -197
rect 563 -216 567 -212
rect 582 -219 586 -190
rect 593 -201 597 -197
rect 593 -216 596 -212
rect 610 -213 613 -209
rect 620 -216 624 -205
rect 640 -213 643 -209
rect 650 -216 654 -205
rect 459 -234 463 -224
rect 470 -231 472 -227
rect 489 -234 493 -224
rect 500 -231 502 -227
rect 459 -237 468 -234
rect 489 -237 498 -234
rect 610 -220 624 -216
rect 640 -220 654 -216
rect 454 -244 478 -240
rect 484 -244 508 -240
rect 560 -243 564 -239
rect 590 -243 594 -239
rect 107 -269 161 -265
rect 167 -269 191 -265
rect 113 -273 117 -269
rect 143 -273 147 -269
rect 173 -273 177 -269
rect 202 -270 256 -266
rect 262 -270 286 -266
rect 112 -324 114 -320
rect -147 -353 -143 -338
rect -136 -346 -133 -342
rect -117 -353 -113 -338
rect 52 -339 54 -335
rect 61 -342 65 -328
rect 82 -339 84 -335
rect 91 -342 95 -328
rect 121 -327 125 -313
rect 142 -324 144 -320
rect 151 -321 155 -313
rect 181 -321 185 -313
rect 208 -274 212 -270
rect 238 -274 242 -270
rect 268 -274 272 -270
rect 151 -325 174 -321
rect 181 -325 190 -321
rect 207 -325 209 -321
rect 151 -327 155 -325
rect 112 -333 114 -329
rect 121 -330 155 -327
rect 181 -328 185 -325
rect 121 -336 125 -330
rect -106 -346 -103 -342
rect 61 -345 95 -342
rect 61 -353 65 -345
rect 91 -353 95 -345
rect -207 -387 -203 -358
rect -196 -369 -192 -365
rect -196 -384 -192 -380
rect -177 -387 -173 -358
rect -166 -369 -162 -365
rect -166 -384 -160 -380
rect -149 -381 -146 -377
rect -139 -384 -135 -373
rect -119 -381 -116 -377
rect -109 -384 -105 -373
rect -149 -388 -135 -384
rect -119 -388 -105 -384
rect -199 -411 -195 -407
rect -169 -411 -165 -407
rect -207 -414 -195 -411
rect -177 -414 -165 -411
rect -242 -421 -218 -417
rect -212 -420 -188 -417
rect -182 -420 -158 -417
rect -152 -420 -128 -417
rect -122 -420 -98 -417
rect -236 -425 -232 -421
rect -228 -473 -224 -465
rect -206 -426 -202 -420
rect -176 -426 -172 -420
rect -146 -426 -142 -420
rect -116 -426 -112 -420
rect -239 -477 -235 -473
rect -228 -477 -219 -473
rect -228 -480 -224 -477
rect -208 -480 -205 -476
rect -198 -487 -194 -466
rect -178 -480 -175 -476
rect -168 -487 -164 -466
rect -148 -480 -145 -476
rect -138 -487 -134 -466
rect -118 -480 -115 -476
rect -108 -487 -104 -466
rect -236 -505 -232 -500
rect -236 -509 -224 -505
rect 216 -328 220 -314
rect 237 -325 239 -321
rect 246 -322 250 -314
rect 276 -322 280 -314
rect 317 -281 321 -250
rect 395 -255 399 -247
rect 429 -255 433 -247
rect 460 -248 464 -244
rect 490 -248 494 -244
rect 552 -246 564 -243
rect 582 -246 594 -243
rect 384 -259 388 -255
rect 395 -259 403 -255
rect 418 -259 422 -255
rect 429 -259 437 -255
rect 328 -263 330 -259
rect 395 -262 399 -259
rect 429 -262 433 -259
rect 328 -272 330 -268
rect 246 -326 269 -322
rect 276 -326 285 -322
rect 246 -328 250 -326
rect 207 -334 209 -330
rect 216 -331 250 -328
rect 276 -329 280 -326
rect 216 -337 220 -331
rect 173 -353 177 -348
rect 173 -357 185 -353
rect 113 -387 117 -376
rect 268 -354 272 -349
rect 268 -358 280 -354
rect 387 -287 391 -282
rect 421 -287 425 -282
rect 387 -291 399 -287
rect 421 -291 433 -287
rect 345 -317 369 -313
rect 351 -321 355 -317
rect 514 -253 538 -249
rect 544 -252 568 -249
rect 574 -252 598 -249
rect 604 -252 628 -249
rect 634 -252 658 -249
rect 520 -257 524 -253
rect 528 -305 532 -297
rect 550 -258 554 -252
rect 580 -258 584 -252
rect 610 -258 614 -252
rect 640 -258 644 -252
rect 664 -253 688 -249
rect 670 -257 674 -253
rect 517 -309 521 -305
rect 528 -309 537 -305
rect 528 -312 532 -309
rect 548 -312 551 -308
rect 459 -339 461 -335
rect 468 -342 472 -328
rect 489 -339 491 -335
rect 498 -342 502 -328
rect 558 -319 562 -298
rect 578 -312 581 -308
rect 588 -319 592 -298
rect 608 -312 611 -308
rect 618 -319 622 -298
rect 638 -312 641 -308
rect 648 -309 652 -298
rect 678 -305 682 -297
rect 664 -309 671 -305
rect 678 -309 687 -305
rect 648 -312 667 -309
rect 678 -312 682 -309
rect 648 -319 652 -312
rect 520 -337 524 -332
rect 520 -341 532 -337
rect 468 -345 502 -342
rect 468 -353 472 -345
rect 498 -353 502 -345
rect 325 -369 329 -361
rect 359 -369 363 -361
rect 325 -373 352 -369
rect 359 -373 368 -369
rect 325 -377 329 -373
rect 359 -376 363 -373
rect 53 -447 57 -433
rect 64 -444 66 -440
rect 83 -447 87 -433
rect 112 -434 114 -430
rect 121 -437 125 -427
rect 208 -388 212 -377
rect 316 -381 318 -377
rect 325 -380 339 -377
rect 325 -384 329 -380
rect 335 -384 339 -380
rect 346 -381 348 -377
rect 317 -408 321 -404
rect 343 -408 347 -404
rect 351 -401 355 -396
rect 351 -405 363 -401
rect 317 -411 347 -408
rect 311 -419 335 -415
rect 325 -423 329 -419
rect 207 -435 209 -431
rect 112 -440 125 -437
rect 216 -438 220 -428
rect 94 -444 96 -440
rect 207 -441 220 -438
rect 107 -447 161 -443
rect 167 -447 191 -443
rect 53 -450 87 -447
rect 53 -460 57 -450
rect 64 -457 66 -453
rect 83 -460 87 -450
rect 113 -451 117 -447
rect 143 -451 147 -447
rect 173 -451 177 -447
rect 203 -448 257 -444
rect 263 -448 287 -444
rect 94 -457 96 -453
rect -146 -522 -142 -507
rect -135 -515 -132 -511
rect -116 -522 -112 -507
rect -105 -515 -102 -511
rect 61 -515 65 -500
rect 91 -515 95 -500
rect 112 -502 114 -498
rect 121 -505 125 -491
rect 142 -502 144 -498
rect 151 -499 155 -491
rect 181 -499 185 -491
rect 209 -452 213 -448
rect 239 -452 243 -448
rect 269 -452 273 -448
rect 151 -503 174 -499
rect 181 -503 190 -499
rect 208 -503 210 -499
rect 151 -505 155 -503
rect 112 -511 114 -507
rect 121 -508 155 -505
rect 181 -506 185 -503
rect 121 -514 125 -508
rect -206 -556 -202 -527
rect -195 -538 -191 -534
rect -195 -553 -191 -549
rect -176 -556 -172 -527
rect -165 -538 -161 -534
rect -165 -553 -159 -549
rect -148 -550 -145 -546
rect -138 -553 -134 -542
rect -118 -550 -115 -546
rect -108 -553 -104 -542
rect -148 -557 -134 -553
rect -118 -557 -104 -553
rect 217 -506 221 -492
rect 238 -503 240 -499
rect 247 -500 251 -492
rect 277 -500 281 -492
rect 247 -504 270 -500
rect 277 -504 286 -500
rect 670 -337 674 -332
rect 610 -354 614 -339
rect 621 -347 624 -343
rect 640 -354 644 -339
rect 670 -341 682 -337
rect 651 -347 654 -343
rect 550 -388 554 -359
rect 561 -370 565 -366
rect 561 -385 565 -381
rect 580 -388 584 -359
rect 591 -370 595 -366
rect 591 -385 594 -381
rect 608 -382 611 -378
rect 618 -385 622 -374
rect 638 -382 641 -378
rect 648 -385 652 -374
rect 608 -389 622 -385
rect 638 -389 652 -385
rect 558 -412 562 -408
rect 588 -412 592 -408
rect 550 -415 562 -412
rect 580 -415 592 -412
rect 514 -421 538 -417
rect 545 -421 569 -418
rect 575 -421 599 -418
rect 605 -421 629 -418
rect 635 -421 659 -418
rect 520 -425 524 -421
rect 460 -447 464 -433
rect 471 -444 473 -440
rect 490 -447 494 -433
rect 501 -444 503 -440
rect 460 -450 494 -447
rect 460 -460 464 -450
rect 471 -457 473 -453
rect 490 -460 494 -450
rect 501 -457 503 -453
rect 528 -473 532 -465
rect 551 -427 555 -421
rect 581 -427 585 -421
rect 611 -427 615 -421
rect 641 -427 645 -421
rect 665 -422 689 -418
rect 671 -426 675 -422
rect 517 -477 521 -473
rect 528 -477 537 -473
rect 528 -480 532 -477
rect 247 -506 251 -504
rect 208 -512 210 -508
rect 217 -509 251 -506
rect 277 -507 281 -504
rect 217 -515 221 -509
rect 173 -531 177 -526
rect 173 -535 185 -531
rect 53 -565 57 -555
rect 64 -562 66 -558
rect 83 -565 87 -555
rect 94 -562 96 -558
rect 113 -565 117 -554
rect 269 -532 273 -527
rect 269 -536 281 -532
rect 317 -534 321 -503
rect 328 -516 330 -512
rect 468 -515 472 -500
rect 498 -515 502 -500
rect 549 -481 552 -477
rect 559 -488 563 -467
rect 579 -481 582 -477
rect 589 -488 593 -467
rect 609 -481 612 -477
rect 619 -488 623 -467
rect 639 -481 642 -477
rect 649 -478 653 -467
rect 679 -474 683 -466
rect 665 -478 672 -474
rect 679 -478 688 -474
rect 649 -481 668 -478
rect 679 -481 683 -478
rect 649 -488 653 -481
rect 520 -505 524 -500
rect 520 -509 532 -505
rect 328 -525 330 -521
rect 53 -568 62 -565
rect 83 -568 92 -565
rect 52 -576 76 -572
rect 82 -576 106 -572
rect -198 -580 -194 -576
rect -168 -580 -164 -576
rect -206 -583 -194 -580
rect -176 -583 -164 -580
rect 58 -580 62 -576
rect 88 -580 92 -576
rect -237 -591 -213 -587
rect -207 -590 -183 -587
rect -177 -590 -153 -587
rect -147 -590 -123 -587
rect -117 -590 -93 -587
rect -231 -595 -227 -591
rect -223 -643 -219 -635
rect -201 -596 -197 -590
rect -171 -596 -167 -590
rect -141 -596 -137 -590
rect -111 -596 -107 -590
rect -234 -647 -230 -643
rect -223 -647 -214 -643
rect -223 -650 -219 -647
rect -203 -650 -200 -646
rect -193 -657 -189 -636
rect -173 -650 -170 -646
rect -163 -657 -159 -636
rect -143 -650 -140 -646
rect -133 -657 -129 -636
rect -113 -650 -110 -646
rect -103 -657 -99 -636
rect -231 -675 -227 -670
rect -231 -679 -219 -675
rect 112 -612 114 -608
rect 121 -615 125 -605
rect 209 -566 213 -555
rect 208 -613 210 -609
rect 112 -618 125 -615
rect 217 -616 221 -606
rect 671 -506 675 -501
rect 611 -523 615 -508
rect 622 -516 625 -512
rect 641 -523 645 -508
rect 671 -510 683 -506
rect 652 -516 655 -512
rect 460 -565 464 -555
rect 471 -562 473 -558
rect 490 -565 494 -555
rect 551 -557 555 -528
rect 562 -539 566 -535
rect 562 -554 566 -550
rect 581 -557 585 -528
rect 592 -539 596 -535
rect 592 -554 595 -550
rect 609 -551 612 -547
rect 619 -554 623 -543
rect 639 -551 642 -547
rect 649 -554 653 -543
rect 501 -562 503 -558
rect 345 -570 369 -566
rect 460 -568 469 -565
rect 490 -568 499 -565
rect 351 -574 355 -570
rect 455 -575 479 -571
rect 485 -575 509 -571
rect 208 -619 221 -616
rect 325 -622 329 -614
rect 359 -622 363 -614
rect 461 -579 465 -575
rect 491 -579 495 -575
rect 609 -558 623 -554
rect 639 -558 653 -554
rect 325 -626 352 -622
rect 359 -626 368 -622
rect 325 -630 329 -626
rect 359 -629 363 -626
rect 316 -634 318 -630
rect 325 -633 339 -630
rect 325 -637 329 -633
rect 57 -671 59 -667
rect 66 -674 70 -660
rect 87 -671 89 -667
rect 96 -674 100 -660
rect 335 -637 339 -633
rect 346 -634 348 -630
rect 317 -661 321 -657
rect 343 -661 347 -657
rect 351 -654 355 -649
rect 351 -658 363 -654
rect 559 -581 563 -577
rect 589 -581 593 -577
rect 551 -584 563 -581
rect 581 -584 593 -581
rect 515 -592 539 -588
rect 550 -591 574 -588
rect 580 -591 604 -588
rect 610 -591 634 -588
rect 640 -591 664 -588
rect 521 -596 525 -592
rect 529 -644 533 -636
rect 556 -597 560 -591
rect 586 -597 590 -591
rect 616 -597 620 -591
rect 646 -597 650 -591
rect 670 -592 694 -588
rect 676 -596 680 -592
rect 518 -648 522 -644
rect 529 -648 538 -644
rect 529 -651 533 -648
rect 554 -651 557 -647
rect 317 -664 347 -661
rect 311 -672 335 -668
rect 460 -670 462 -666
rect 66 -677 100 -674
rect 325 -676 329 -672
rect -141 -692 -137 -677
rect -130 -685 -127 -681
rect -111 -692 -107 -677
rect -100 -685 -97 -681
rect 66 -685 70 -677
rect 96 -685 100 -677
rect -201 -726 -197 -697
rect -190 -708 -186 -704
rect -190 -723 -186 -719
rect -171 -726 -167 -697
rect -160 -708 -156 -704
rect -160 -723 -154 -719
rect -143 -720 -140 -716
rect -133 -723 -129 -712
rect -113 -720 -110 -716
rect -103 -723 -99 -712
rect -143 -727 -129 -723
rect -113 -727 -99 -723
rect -193 -750 -189 -746
rect -163 -750 -159 -746
rect -201 -753 -189 -750
rect -171 -753 -159 -750
rect -234 -762 -210 -758
rect -204 -761 -180 -758
rect -174 -761 -150 -758
rect -144 -761 -120 -758
rect -114 -761 -90 -758
rect -228 -766 -224 -762
rect -220 -814 -216 -806
rect -198 -767 -194 -761
rect -168 -767 -164 -761
rect -138 -767 -134 -761
rect -108 -767 -104 -761
rect 469 -673 473 -659
rect 490 -670 492 -666
rect 499 -673 503 -659
rect 469 -676 503 -673
rect 469 -684 473 -676
rect 499 -684 503 -676
rect 564 -658 568 -637
rect 584 -651 587 -647
rect 594 -658 598 -637
rect 614 -651 617 -647
rect 624 -658 628 -637
rect 644 -651 647 -647
rect 654 -648 658 -637
rect 684 -644 688 -636
rect 670 -648 677 -644
rect 684 -648 693 -644
rect 654 -651 673 -648
rect 684 -651 688 -648
rect 654 -658 658 -651
rect 521 -676 525 -671
rect 521 -680 533 -676
rect -231 -818 -227 -814
rect -220 -818 -211 -814
rect -220 -821 -216 -818
rect -200 -821 -197 -817
rect -190 -828 -186 -807
rect -170 -821 -167 -817
rect -160 -828 -156 -807
rect -140 -821 -137 -817
rect -130 -828 -126 -807
rect -110 -821 -107 -817
rect -100 -828 -96 -807
rect -228 -846 -224 -841
rect -228 -850 -216 -846
rect 58 -779 62 -765
rect 69 -776 71 -772
rect 88 -779 92 -765
rect 99 -776 101 -772
rect 58 -782 92 -779
rect 58 -792 62 -782
rect 69 -789 71 -785
rect 88 -792 92 -782
rect 99 -789 101 -785
rect 317 -787 321 -756
rect 676 -676 680 -671
rect 616 -693 620 -678
rect 627 -686 630 -682
rect 646 -693 650 -678
rect 676 -680 688 -676
rect 657 -686 660 -682
rect 556 -727 560 -698
rect 567 -709 571 -705
rect 567 -724 571 -720
rect 586 -727 590 -698
rect 597 -709 601 -705
rect 597 -724 600 -720
rect 614 -721 617 -717
rect 624 -724 628 -713
rect 644 -721 647 -717
rect 654 -724 658 -713
rect 614 -728 628 -724
rect 644 -728 658 -724
rect 564 -751 568 -747
rect 594 -751 598 -747
rect 556 -754 568 -751
rect 586 -754 598 -751
rect 328 -769 330 -765
rect 328 -778 330 -774
rect 461 -778 465 -764
rect 472 -775 474 -771
rect 491 -778 495 -764
rect 502 -775 504 -771
rect 461 -781 495 -778
rect 66 -847 70 -832
rect 96 -847 100 -832
rect -138 -863 -134 -848
rect -127 -856 -124 -852
rect -108 -863 -104 -848
rect -97 -856 -94 -852
rect -198 -897 -194 -868
rect -187 -879 -183 -875
rect -187 -894 -183 -890
rect -168 -897 -164 -868
rect -157 -879 -153 -875
rect -157 -894 -151 -890
rect -140 -891 -137 -887
rect -130 -894 -126 -883
rect -110 -891 -107 -887
rect -100 -894 -96 -883
rect -140 -898 -126 -894
rect -110 -898 -96 -894
rect 461 -791 465 -781
rect 472 -788 474 -784
rect 491 -791 495 -781
rect 502 -788 504 -784
rect 345 -823 369 -819
rect 351 -827 355 -823
rect 469 -846 473 -831
rect 499 -846 503 -831
rect 325 -875 329 -867
rect 359 -875 363 -867
rect 325 -879 352 -875
rect 359 -879 368 -875
rect 325 -883 329 -879
rect 359 -882 363 -879
rect 316 -887 318 -883
rect 325 -886 339 -883
rect 58 -897 62 -887
rect 69 -894 71 -890
rect 88 -897 92 -887
rect 325 -890 329 -886
rect 99 -894 101 -890
rect 58 -900 67 -897
rect 88 -900 97 -897
rect 56 -909 80 -905
rect 86 -909 110 -905
rect -190 -921 -186 -917
rect -160 -921 -156 -917
rect -198 -924 -186 -921
rect -168 -924 -156 -921
rect 62 -913 66 -909
rect 92 -913 96 -909
rect 335 -890 339 -886
rect 346 -887 348 -883
rect -232 -933 -208 -929
rect -202 -932 -178 -929
rect -172 -932 -148 -929
rect -142 -932 -118 -929
rect -112 -932 -88 -929
rect -226 -937 -222 -933
rect -218 -985 -214 -977
rect -196 -938 -192 -932
rect -166 -938 -162 -932
rect -136 -938 -132 -932
rect -106 -938 -102 -932
rect -229 -989 -225 -985
rect -218 -989 -209 -985
rect -218 -992 -214 -989
rect -198 -992 -195 -988
rect -188 -999 -184 -978
rect -168 -992 -165 -988
rect -158 -999 -154 -978
rect -138 -992 -135 -988
rect -128 -999 -124 -978
rect -108 -992 -105 -988
rect -98 -999 -94 -978
rect 317 -914 321 -910
rect 343 -914 347 -910
rect 461 -896 465 -886
rect 472 -893 474 -889
rect 491 -896 495 -886
rect 502 -893 504 -889
rect 461 -899 470 -896
rect 491 -899 500 -896
rect 351 -907 355 -902
rect 454 -906 478 -902
rect 484 -906 508 -902
rect 351 -911 363 -907
rect 460 -910 464 -906
rect 490 -910 494 -906
rect 317 -917 347 -914
rect -226 -1017 -222 -1012
rect -226 -1021 -214 -1017
rect 61 -1004 63 -1000
rect 70 -1007 74 -993
rect 91 -1004 93 -1000
rect 100 -1007 104 -993
rect 459 -1001 461 -997
rect 70 -1010 104 -1007
rect 70 -1018 74 -1010
rect 100 -1018 104 -1010
rect 468 -1004 472 -990
rect 489 -1001 491 -997
rect 498 -1004 502 -990
rect 468 -1007 502 -1004
rect 468 -1015 472 -1007
rect 498 -1015 502 -1007
rect -136 -1034 -132 -1019
rect -125 -1027 -122 -1023
rect -106 -1034 -102 -1019
rect -95 -1027 -92 -1023
rect -196 -1068 -192 -1039
rect -185 -1050 -181 -1046
rect -185 -1065 -181 -1061
rect -166 -1068 -162 -1039
rect -155 -1050 -151 -1046
rect -155 -1065 -149 -1061
rect -138 -1062 -135 -1058
rect -128 -1065 -124 -1054
rect -108 -1062 -105 -1058
rect -98 -1065 -94 -1054
rect -138 -1069 -124 -1065
rect -108 -1069 -94 -1065
rect -188 -1092 -184 -1088
rect -158 -1092 -154 -1088
rect -196 -1095 -184 -1092
rect -166 -1095 -154 -1092
rect -229 -1105 -205 -1101
rect -199 -1104 -175 -1101
rect -169 -1104 -145 -1101
rect -139 -1104 -115 -1101
rect -109 -1104 -85 -1101
rect -223 -1109 -219 -1105
rect -215 -1157 -211 -1149
rect -193 -1110 -189 -1104
rect -163 -1110 -159 -1104
rect -133 -1110 -129 -1104
rect -103 -1110 -99 -1104
rect -226 -1161 -222 -1157
rect -215 -1161 -206 -1157
rect -215 -1164 -211 -1161
rect -195 -1164 -192 -1160
rect -185 -1171 -181 -1150
rect -165 -1164 -162 -1160
rect -155 -1171 -151 -1150
rect -135 -1164 -132 -1160
rect -125 -1171 -121 -1150
rect -105 -1164 -102 -1160
rect -95 -1171 -91 -1150
rect 62 -1112 66 -1098
rect 73 -1109 75 -1105
rect 92 -1112 96 -1098
rect 103 -1109 105 -1105
rect 460 -1109 464 -1095
rect 471 -1106 473 -1102
rect 490 -1109 494 -1095
rect 501 -1106 503 -1102
rect 62 -1115 96 -1112
rect 62 -1125 66 -1115
rect 73 -1122 75 -1118
rect 92 -1125 96 -1115
rect 460 -1112 494 -1109
rect 103 -1122 105 -1118
rect 460 -1122 464 -1112
rect 471 -1119 473 -1115
rect 490 -1122 494 -1112
rect 501 -1119 503 -1115
rect -223 -1189 -219 -1184
rect -223 -1193 -211 -1189
rect 70 -1180 74 -1165
rect 100 -1180 104 -1165
rect 468 -1177 472 -1162
rect 498 -1177 502 -1162
rect -133 -1206 -129 -1191
rect -122 -1199 -119 -1195
rect -103 -1206 -99 -1191
rect -92 -1199 -89 -1195
rect -193 -1240 -189 -1211
rect -182 -1222 -178 -1218
rect -182 -1237 -178 -1233
rect -163 -1240 -159 -1211
rect -152 -1222 -148 -1218
rect -152 -1237 -146 -1233
rect -135 -1234 -132 -1230
rect -125 -1237 -121 -1226
rect -105 -1234 -102 -1230
rect -95 -1237 -91 -1226
rect 62 -1230 66 -1220
rect 73 -1227 75 -1223
rect 92 -1230 96 -1220
rect 103 -1227 105 -1223
rect 460 -1227 464 -1217
rect 471 -1224 473 -1220
rect 490 -1227 494 -1217
rect 501 -1224 503 -1220
rect 460 -1230 469 -1227
rect 490 -1230 499 -1227
rect 62 -1233 71 -1230
rect 92 -1233 101 -1230
rect -135 -1241 -121 -1237
rect -105 -1241 -91 -1237
rect -185 -1264 -181 -1260
rect -155 -1264 -151 -1260
rect -193 -1267 -181 -1264
rect -163 -1267 -151 -1264
<< labels >>
rlabel metal1 -19 1 -19 1 1 gnd
rlabel metal1 -14 -96 -14 -96 1 gnd
rlabel metal1 15 1 15 1 1 gnd
rlabel metal1 20 -96 20 -96 1 gnd
rlabel metal1 -13 -192 -13 -192 1 gnd
rlabel metal1 -8 -289 -8 -289 1 gnd
rlabel metal1 21 -192 21 -192 1 gnd
rlabel metal1 26 -289 26 -289 1 gnd
rlabel metal1 -25 33 -25 33 1 A0
rlabel metal1 -8 33 -8 33 1 A0_n
rlabel metal1 10 33 10 33 1 B0
rlabel metal1 26 33 26 33 1 B0_n
rlabel metal1 -19 -64 -19 -64 1 A1
rlabel metal1 -5 -64 -5 -64 1 A1_n
rlabel metal1 31 -64 31 -64 1 B1_n
rlabel metal1 15 -64 15 -64 1 B1
rlabel metal1 -18 -160 -18 -160 1 A2
rlabel metal1 -2 -160 -2 -160 1 A2_n
rlabel metal1 16 -160 16 -160 1 B2
rlabel metal1 31 -160 31 -160 1 B2_n
rlabel metal1 -13 -257 -13 -257 1 A3
rlabel metal1 2 -257 2 -257 1 A3_n
rlabel metal1 20 -257 20 -257 1 B3
rlabel metal1 36 -257 36 -257 7 B3_n
rlabel metal1 -22 90 -22 90 5 vdd
rlabel metal1 12 90 12 90 5 vdd
rlabel metal1 50 90 50 90 5 vdd
rlabel metal1 79 90 79 90 5 vdd
rlabel metal1 -16 -103 -16 -103 5 vdd
rlabel metal1 18 -103 18 -103 5 vdd
rlabel metal1 -11 -200 -11 -200 5 vdd
rlabel metal1 23 -200 23 -200 5 vdd
rlabel metal1 -17 -7 -17 -7 5 vdd
rlabel metal1 17 -7 17 -7 5 vdd
rlabel metal1 52 -235 52 -235 1 gnd
rlabel metal1 82 -235 82 -235 1 gnd
rlabel metal1 54 -241 54 -241 5 vdd
rlabel metal1 83 -241 83 -241 5 vdd
rlabel metal1 56 -566 56 -566 1 gnd
rlabel metal1 86 -566 86 -566 1 gnd
rlabel metal1 59 -573 59 -573 5 vdd
rlabel metal1 88 -573 88 -573 5 vdd
rlabel metal1 61 -898 61 -898 1 gnd
rlabel metal1 91 -898 91 -898 1 gnd
rlabel metal1 63 -906 63 -906 5 vdd
rlabel metal1 92 -906 92 -906 5 vdd
rlabel metal1 65 -1231 65 -1231 1 gnd
rlabel metal1 95 -1231 95 -1231 1 gnd
rlabel metal1 49 -6 49 -6 1 A0
rlabel metal1 79 -6 79 -6 1 B0
rlabel metal1 61 -111 61 -111 1 A0_n
rlabel metal1 91 -111 91 -111 1 B0_n
rlabel metal1 61 -124 61 -124 1 A0
rlabel metal1 91 -124 91 -124 1 A0_n
rlabel metal1 61 -229 61 -229 1 B0
rlabel metal1 91 -229 91 -229 1 B0_n
rlabel metal1 53 -338 53 -338 1 A1
rlabel metal1 83 -337 83 -337 1 B1
rlabel metal1 65 -442 65 -442 1 A1_n
rlabel metal1 95 -442 95 -442 1 B1_n
rlabel metal1 65 -455 65 -455 1 A1
rlabel metal1 95 -454 95 -454 1 A1_n
rlabel metal1 65 -560 65 -560 1 B1
rlabel metal1 95 -560 95 -560 1 B1_n
rlabel metal1 58 -669 58 -669 1 A2
rlabel metal1 88 -669 88 -669 1 B2
rlabel metal1 70 -775 70 -775 1 A2_n
rlabel metal1 100 -774 100 -774 1 B2_n
rlabel metal1 90 -781 90 -781 1 P2
rlabel metal1 70 -788 70 -788 1 A2
rlabel metal1 100 -786 100 -786 1 A2_n
rlabel metal1 70 -892 70 -892 1 B2
rlabel metal1 100 -892 100 -892 1 B2_n
rlabel metal1 62 -1003 62 -1003 1 A3
rlabel metal1 92 -1003 92 -1003 1 B3
rlabel metal1 74 -1107 74 -1107 1 A3_n
rlabel metal1 104 -1107 104 -1107 1 B3_n
rlabel metal1 94 -1114 94 -1114 1 P3
rlabel metal1 74 -1120 74 -1120 1 A3
rlabel metal1 104 -1120 104 -1120 1 A3_n
rlabel metal1 74 -1225 74 -1225 1 B3
rlabel metal1 104 -1225 104 -1225 1 B3_n
rlabel metal1 85 -448 85 -448 1 P1
rlabel metal1 81 -117 81 -117 1 P0
rlabel metal1 116 -82 116 -82 1 gnd
rlabel metal1 128 -88 128 -88 5 vdd
rlabel metal1 116 -260 116 -260 1 gnd
rlabel metal1 132 -266 132 -266 5 vdd
rlabel metal1 120 -438 120 -438 1 gnd
rlabel metal1 132 -444 132 -444 5 vdd
rlabel metal1 120 -616 120 -616 1 gnd
rlabel metal1 173 1 173 1 1 gnd
rlabel metal1 170 90 170 90 5 vdd
rlabel metal1 128 90 128 90 5 vdd
rlabel metal1 173 -177 173 -177 1 gnd
rlabel metal1 170 -88 170 -88 5 vdd
rlabel metal1 177 -355 177 -355 1 gnd
rlabel metal1 174 -266 174 -266 5 vdd
rlabel metal1 177 -533 177 -533 1 gnd
rlabel metal1 174 -444 174 -444 5 vdd
rlabel metal1 109 34 109 34 1 A0
rlabel metal1 139 34 139 34 1 B0
rlabel metal1 109 25 109 25 1 A0
rlabel metal1 109 -76 109 -76 1 B0
rlabel metal1 185 33 185 33 1 G0
rlabel metal1 109 -144 109 -144 1 A1
rlabel metal1 139 -144 139 -144 1 B1
rlabel metal1 109 -153 109 -153 1 A1
rlabel metal1 184 -145 184 -145 1 G1
rlabel metal1 109 -254 109 -254 1 B1
rlabel metal1 113 -322 113 -322 1 A2
rlabel metal1 143 -322 143 -322 1 B2
rlabel metal1 113 -331 113 -331 1 A2
rlabel metal1 188 -323 188 -323 7 G2
rlabel metal1 113 -432 113 -432 1 B2
rlabel metal1 113 -500 113 -500 1 A3
rlabel metal1 143 -500 143 -500 1 B3
rlabel metal1 113 -509 113 -509 1 A3
rlabel metal1 188 -501 188 -501 7 G3
rlabel metal1 113 -610 113 -610 1 B3
rlabel metal1 218 -82 218 -82 1 gnd
rlabel metal1 275 1 275 1 1 gnd
rlabel metal1 272 90 272 90 5 vdd
rlabel metal1 230 90 230 90 5 vdd
rlabel metal1 276 -177 276 -177 1 gnd
rlabel metal1 273 -88 273 -88 5 vdd
rlabel metal1 231 -88 231 -88 5 vdd
rlabel metal1 215 -439 215 -439 1 gnd
rlabel metal1 272 -356 272 -356 1 gnd
rlabel metal1 269 -267 269 -267 5 vdd
rlabel metal1 227 -267 227 -267 5 vdd
rlabel metal1 216 -617 216 -617 1 gnd
rlabel metal1 273 -534 273 -534 1 gnd
rlabel metal1 270 -445 270 -445 5 vdd
rlabel metal1 228 -445 228 -445 5 vdd
rlabel metal1 218 -261 218 -261 1 gnd
rlabel metal1 211 34 211 34 1 P0
rlabel metal1 211 25 211 25 1 P0
rlabel metal1 241 34 241 34 1 gnd
rlabel metal1 211 -76 211 -76 1 gnd
rlabel metal1 287 33 287 33 7 PC0
rlabel metal1 212 -144 212 -144 1 P1
rlabel metal1 212 -153 212 -153 1 P1
rlabel metal1 242 -144 242 -144 1 C1
rlabel metal1 212 -254 212 -254 1 C1
rlabel metal1 208 -323 208 -323 1 P2
rlabel metal1 208 -332 208 -332 1 P2
rlabel metal1 238 -323 238 -323 1 C2
rlabel metal1 208 -433 208 -433 1 C2
rlabel metal1 287 -145 287 -145 7 PC1
rlabel metal1 283 -325 283 -325 1 PC2
rlabel metal1 209 -501 209 -501 1 P3
rlabel metal1 209 -510 209 -510 1 P3
rlabel metal1 239 -501 239 -501 1 C3
rlabel metal1 285 -502 285 -502 7 PC3
rlabel metal1 331 -156 331 -156 1 gnd
rlabel metal1 323 90 323 90 5 vdd
rlabel metal1 331 -409 331 -409 1 gnd
rlabel metal1 323 -163 323 -163 5 vdd
rlabel metal1 331 -662 331 -662 1 gnd
rlabel metal1 323 -416 323 -416 5 vdd
rlabel metal1 331 -915 331 -915 1 gnd
rlabel metal1 323 -669 323 -669 5 vdd
rlabel metal1 355 -149 355 -149 1 gnd
rlabel metal1 352 -60 352 -60 5 vdd
rlabel metal1 355 -403 355 -403 1 gnd
rlabel metal1 352 -314 352 -314 5 vdd
rlabel metal1 355 -656 355 -656 1 gnd
rlabel metal1 352 -567 352 -567 5 vdd
rlabel metal1 355 -909 355 -909 1 gnd
rlabel metal1 352 -820 352 -820 5 vdd
rlabel metal1 329 -8 329 -8 1 PC0
rlabel metal1 329 -17 329 -17 1 G0
rlabel metal1 317 -127 317 -127 1 PC0
rlabel metal1 347 -126 347 -126 1 G0
rlabel metal1 366 -117 366 -117 7 C1
rlabel metal1 329 -261 329 -261 1 PC1
rlabel metal1 329 -270 329 -270 1 G1
rlabel metal1 317 -379 317 -379 1 PC1
rlabel metal1 347 -379 347 -379 1 G1
rlabel metal1 366 -371 366 -371 7 C2
rlabel metal1 329 -514 329 -514 1 PC2
rlabel metal1 329 -523 329 -523 1 G2
rlabel metal1 317 -632 317 -632 1 PC2
rlabel metal1 347 -632 347 -632 1 G2
rlabel metal1 366 -624 366 -624 7 C3
rlabel metal1 329 -767 329 -767 1 PC3
rlabel metal1 329 -776 329 -776 1 G3
rlabel metal1 317 -885 317 -885 1 PC3
rlabel metal1 347 -885 347 -885 1 G3
rlabel metal1 380 1 380 1 1 gnd
rlabel metal1 385 -96 385 -96 1 gnd
rlabel metal1 414 1 414 1 1 gnd
rlabel metal1 419 -96 419 -96 1 gnd
rlabel metal1 386 -192 386 -192 1 gnd
rlabel metal1 391 -289 391 -289 1 gnd
rlabel metal1 420 -192 420 -192 1 gnd
rlabel metal1 425 -289 425 -289 1 gnd
rlabel metal1 377 90 377 90 5 vdd
rlabel metal1 411 90 411 90 5 vdd
rlabel metal1 383 -103 383 -103 5 vdd
rlabel metal1 417 -103 417 -103 5 vdd
rlabel metal1 388 -200 388 -200 5 vdd
rlabel metal1 422 -200 422 -200 5 vdd
rlabel metal1 382 -7 382 -7 5 vdd
rlabel metal1 416 -7 416 -7 5 vdd
rlabel metal1 374 33 374 33 1 P0
rlabel metal1 391 33 391 33 1 P0_n
rlabel metal1 409 33 409 33 1 gnd
rlabel metal1 425 33 425 33 1 C0_n
rlabel metal1 380 -64 380 -64 1 P1
rlabel metal1 394 -64 394 -64 1 P1_n
rlabel metal1 414 -64 414 -64 1 C1
rlabel metal1 430 -64 430 -64 1 C1_n
rlabel metal1 381 -160 381 -160 1 P2
rlabel metal1 397 -160 397 -160 1 P2_n
rlabel metal1 415 -160 415 -160 1 C2
rlabel metal1 430 -160 430 -160 1 C2_n
rlabel metal1 386 -257 386 -257 1 P3
rlabel metal1 401 -257 401 -257 1 P3_n
rlabel metal1 419 -257 419 -257 1 C3
rlabel metal1 435 -257 435 -257 7 C3_n
rlabel metal1 460 90 460 90 5 vdd
rlabel metal1 489 90 489 90 5 vdd
rlabel metal1 462 -235 462 -235 1 gnd
rlabel metal1 492 -235 492 -235 1 gnd
rlabel metal1 461 -241 461 -241 5 vdd
rlabel metal1 490 -241 490 -241 5 vdd
rlabel metal1 463 -566 463 -566 1 gnd
rlabel metal1 493 -566 493 -566 1 gnd
rlabel metal1 462 -572 462 -572 5 vdd
rlabel metal1 491 -572 491 -572 5 vdd
rlabel metal1 464 -897 464 -897 1 gnd
rlabel metal1 494 -897 494 -897 1 gnd
rlabel metal1 461 -903 461 -903 5 vdd
rlabel metal1 490 -903 490 -903 5 vdd
rlabel metal1 463 -1228 463 -1228 1 gnd
rlabel metal1 493 -1228 493 -1228 1 gnd
rlabel metal1 459 -6 459 -6 1 P0
rlabel metal1 489 -6 489 -6 1 gnd
rlabel metal1 471 -111 471 -111 1 P0_n
rlabel metal1 501 -111 501 -111 1 C0_n
rlabel metal1 501 -124 501 -124 1 P0_n
rlabel metal1 471 -124 471 -124 1 P0
rlabel metal1 491 -117 491 -117 1 Sum0_unlatched
rlabel metal1 471 -229 471 -229 1 gnd
rlabel metal1 501 -229 501 -229 1 C0_n
rlabel metal1 460 -337 460 -337 1 P1
rlabel metal1 490 -337 490 -337 1 C1
rlabel metal1 472 -442 472 -442 1 P1_n
rlabel metal1 502 -442 502 -442 1 C1_n
rlabel metal1 492 -448 492 -448 1 Sum1_unlatched
rlabel metal1 472 -455 472 -455 1 P1
rlabel metal1 502 -455 502 -455 1 P1_n
rlabel metal1 472 -560 472 -560 1 C1
rlabel metal1 502 -560 502 -560 1 C1_n
rlabel metal1 461 -668 461 -668 1 P2
rlabel metal1 491 -668 491 -668 1 C2
rlabel metal1 473 -773 473 -773 1 P2_n
rlabel metal1 503 -773 503 -773 1 C2_n
rlabel metal1 503 -786 503 -786 1 P2_n
rlabel metal1 473 -786 473 -786 1 P2
rlabel metal1 493 -779 493 -779 1 Sum2_unlatched
rlabel metal1 366 -877 366 -877 1 Cout_unlatched
rlabel metal1 473 -891 473 -891 1 C2
rlabel metal1 503 -891 503 -891 1 C2_n
rlabel metal1 460 -999 460 -999 1 P3
rlabel metal1 490 -999 490 -999 1 C3
rlabel metal1 472 -1104 472 -1104 1 P3_n
rlabel metal1 502 -1104 502 -1104 1 C3_n
rlabel metal1 472 -1117 472 -1117 1 P3
rlabel metal1 502 -1117 502 -1117 1 P3_n
rlabel metal1 472 -1222 472 -1222 1 C3
rlabel metal1 502 -1222 502 -1222 1 C3_n
rlabel metal1 492 -1110 492 -1110 1 Sum3_unlatched
rlabel metal1 209 -611 209 -611 1 C3
rlabel metal1 -84 2 -84 2 1 gnd
rlabel metal1 -79 -95 -79 -95 1 gnd
rlabel metal1 -50 2 -50 2 1 gnd
rlabel metal1 -45 -95 -45 -95 1 gnd
rlabel metal1 -78 -191 -78 -191 1 gnd
rlabel metal1 -73 -288 -73 -288 1 gnd
rlabel metal1 -44 -191 -44 -191 1 gnd
rlabel metal1 -39 -288 -39 -288 1 gnd
rlabel metal1 -87 91 -87 91 5 vdd
rlabel metal1 -53 91 -53 91 5 vdd
rlabel metal1 -81 -102 -81 -102 5 vdd
rlabel metal1 -47 -102 -47 -102 5 vdd
rlabel metal1 -76 -199 -76 -199 5 vdd
rlabel metal1 -42 -199 -42 -199 5 vdd
rlabel metal1 -82 -6 -82 -6 5 vdd
rlabel metal1 -48 -6 -48 -6 5 vdd
rlabel metal1 -195 -27 -195 -27 1 CLK
rlabel metal1 -204 90 -204 90 1 vdd
rlabel metal1 -165 -27 -165 -27 1 CLK
rlabel metal1 -174 90 -174 90 1 vdd
rlabel metal1 -198 -73 -198 -73 1 gnd
rlabel metal1 -168 -73 -168 -73 1 gnd
rlabel metal1 -136 -4 -136 -4 1 CLK
rlabel metal1 -143 -46 -143 -46 1 gnd
rlabel metal1 -149 91 -149 91 1 vdd
rlabel metal1 -106 -4 -106 -4 1 CLK
rlabel metal1 -113 -46 -113 -46 1 gnd
rlabel metal1 -119 91 -119 91 1 vdd
rlabel metal1 -192 -198 -192 -198 1 CLK
rlabel metal1 -201 -81 -201 -81 1 vdd
rlabel metal1 -162 -198 -162 -198 1 CLK
rlabel metal1 -171 -81 -171 -81 1 vdd
rlabel metal1 -195 -244 -195 -244 1 gnd
rlabel metal1 -165 -244 -165 -244 1 gnd
rlabel metal1 -133 -175 -133 -175 1 CLK
rlabel metal1 -140 -217 -140 -217 1 gnd
rlabel metal1 -146 -80 -146 -80 1 vdd
rlabel metal1 -103 -175 -103 -175 1 CLK
rlabel metal1 -110 -217 -110 -217 1 gnd
rlabel metal1 -116 -80 -116 -80 1 vdd
rlabel metal1 -194 -367 -194 -367 1 CLK
rlabel metal1 -203 -250 -203 -250 1 vdd
rlabel metal1 -164 -367 -164 -367 1 CLK
rlabel metal1 -173 -250 -173 -250 1 vdd
rlabel metal1 -197 -413 -197 -413 1 gnd
rlabel metal1 -167 -413 -167 -413 1 gnd
rlabel metal1 -135 -344 -135 -344 1 CLK
rlabel metal1 -142 -386 -142 -386 1 gnd
rlabel metal1 -148 -249 -148 -249 1 vdd
rlabel metal1 -105 -344 -105 -344 1 CLK
rlabel metal1 -112 -386 -112 -386 1 gnd
rlabel metal1 -118 -249 -118 -249 1 vdd
rlabel metal1 -193 -536 -193 -536 1 CLK
rlabel metal1 -202 -419 -202 -419 1 vdd
rlabel metal1 -163 -536 -163 -536 1 CLK
rlabel metal1 -172 -419 -172 -419 1 vdd
rlabel metal1 -196 -582 -196 -582 1 gnd
rlabel metal1 -166 -582 -166 -582 1 gnd
rlabel metal1 -134 -513 -134 -513 1 CLK
rlabel metal1 -141 -555 -141 -555 1 gnd
rlabel metal1 -147 -418 -147 -418 1 vdd
rlabel metal1 -104 -513 -104 -513 1 CLK
rlabel metal1 -111 -555 -111 -555 1 gnd
rlabel metal1 -117 -418 -117 -418 1 vdd
rlabel metal1 -188 -706 -188 -706 1 CLK
rlabel metal1 -197 -589 -197 -589 1 vdd
rlabel metal1 -158 -706 -158 -706 1 CLK
rlabel metal1 -167 -589 -167 -589 1 vdd
rlabel metal1 -191 -752 -191 -752 1 gnd
rlabel metal1 -161 -752 -161 -752 1 gnd
rlabel metal1 -129 -683 -129 -683 1 CLK
rlabel metal1 -136 -725 -136 -725 1 gnd
rlabel metal1 -142 -588 -142 -588 1 vdd
rlabel metal1 -99 -683 -99 -683 1 CLK
rlabel metal1 -106 -725 -106 -725 1 gnd
rlabel metal1 -112 -588 -112 -588 1 vdd
rlabel metal1 -206 -140 -206 -140 1 B0_unlatched
rlabel metal1 -203 -206 -203 -206 1 Bb0
rlabel metal1 -163 -213 -163 -213 1 Bb0
rlabel metal1 -176 -140 -176 -140 1 Bb0
rlabel metal1 -146 -210 -146 -210 1 Dnb0
rlabel metal1 -145 -140 -145 -140 1 Dnb0
rlabel metal1 -135 -142 -135 -142 1 Ab0
rlabel metal1 -116 -140 -116 -140 1 Ab0
rlabel metal1 -116 -210 -116 -210 1 Ab0
rlabel metal1 -209 31 -209 31 3 A0_unlatched
rlabel metal1 -206 -35 -206 -35 1 Ba0
rlabel metal1 -166 -42 -166 -42 1 Ba0
rlabel metal1 -179 31 -179 31 1 Ba0
rlabel metal1 -148 31 -148 31 1 Dna0
rlabel metal1 -149 -39 -149 -39 1 Dna0
rlabel metal1 -138 29 -138 29 1 Aa0
rlabel metal1 -119 31 -119 31 1 Aa0
rlabel metal1 -119 -39 -119 -39 1 Aa0
rlabel metal1 -208 -309 -208 -309 1 A1_unlatched
rlabel metal1 -194 -42 -194 -42 1 A0_unlatched
rlabel metal1 -193 -382 -193 -382 1 A1_unlatched
rlabel metal1 -205 -375 -205 -375 1 Ba1
rlabel metal1 -165 -382 -165 -382 1 Ba1
rlabel metal1 -178 -309 -178 -309 1 Ba1
rlabel metal1 -147 -309 -147 -309 1 Dna1
rlabel metal1 -148 -379 -148 -379 1 Dna1
rlabel metal1 -137 -311 -137 -311 1 Aa1
rlabel metal1 -118 -309 -118 -309 1 Aa1
rlabel metal1 -118 -379 -118 -379 1 Aa1
rlabel metal1 -117 -478 -117 -478 1 Ab1
rlabel metal1 -117 -548 -117 -548 1 Ab1
rlabel metal1 -136 -480 -136 -480 1 Ab1
rlabel metal1 -146 -478 -146 -478 1 Dnb1
rlabel metal1 -147 -548 -147 -548 1 Dnb1
rlabel metal1 -164 -551 -164 -551 1 Bb1
rlabel metal1 -177 -478 -177 -478 1 Bb1
rlabel metal1 -207 -478 -207 -478 1 B1_unlatched
rlabel metal1 -192 -551 -192 -551 1 B1_unlatched
rlabel metal1 -204 -544 -204 -544 1 Bb1
rlabel metal1 -202 -648 -202 -648 1 A2_unlatched
rlabel metal1 -199 -714 -199 -714 1 Ba2
rlabel metal1 -187 -721 -187 -721 1 A2_unlatched
rlabel metal1 -159 -721 -159 -721 1 Ba2
rlabel metal1 -172 -648 -172 -648 1 Ba2
rlabel metal1 -141 -648 -141 -648 1 Dna2
rlabel metal1 -131 -650 -131 -650 1 Aa2
rlabel metal1 -142 -718 -142 -718 1 Dna2
rlabel metal1 -112 -718 -112 -718 1 Aa2
rlabel metal1 -112 -648 -112 -648 1 Aa2
rlabel metal1 -185 -877 -185 -877 1 CLK
rlabel metal1 -194 -760 -194 -760 1 vdd
rlabel metal1 -155 -877 -155 -877 1 CLK
rlabel metal1 -164 -760 -164 -760 1 vdd
rlabel metal1 -188 -923 -188 -923 1 gnd
rlabel metal1 -158 -923 -158 -923 1 gnd
rlabel metal1 -126 -854 -126 -854 1 CLK
rlabel metal1 -133 -896 -133 -896 1 gnd
rlabel metal1 -139 -759 -139 -759 1 vdd
rlabel metal1 -96 -854 -96 -854 1 CLK
rlabel metal1 -103 -896 -103 -896 1 gnd
rlabel metal1 -109 -759 -109 -759 1 vdd
rlabel metal1 -199 -819 -199 -819 1 B2_unlatched
rlabel metal1 -184 -892 -184 -892 1 B2_unlatched
rlabel metal1 -196 -885 -196 -885 1 Bb2
rlabel metal1 -156 -892 -156 -892 1 Bb2
rlabel metal1 -169 -819 -169 -819 1 Bb2
rlabel metal1 -138 -819 -138 -819 1 Dnb2
rlabel metal1 -128 -821 -128 -821 1 Ab2
rlabel metal1 -139 -889 -139 -889 1 Dnb2
rlabel metal1 -109 -889 -109 -889 1 Ab2
rlabel metal1 -109 -819 -109 -819 1 Ab2
rlabel metal1 -183 -1048 -183 -1048 1 CLK
rlabel metal1 -192 -931 -192 -931 1 vdd
rlabel metal1 -153 -1048 -153 -1048 1 CLK
rlabel metal1 -162 -931 -162 -931 1 vdd
rlabel metal1 -186 -1094 -186 -1094 1 gnd
rlabel metal1 -156 -1094 -156 -1094 1 gnd
rlabel metal1 -124 -1025 -124 -1025 1 CLK
rlabel metal1 -131 -1067 -131 -1067 1 gnd
rlabel metal1 -137 -930 -137 -930 1 vdd
rlabel metal1 -94 -1025 -94 -1025 1 CLK
rlabel metal1 -101 -1067 -101 -1067 1 gnd
rlabel metal1 -107 -930 -107 -930 1 vdd
rlabel metal1 -197 -990 -197 -990 1 A3_unlatched
rlabel metal1 -194 -1056 -194 -1056 1 Ba3
rlabel metal1 -182 -1063 -182 -1063 1 A3_unlatched
rlabel metal1 -154 -1063 -154 -1063 1 Ba3
rlabel metal1 -167 -990 -167 -990 1 Ba3
rlabel metal1 -136 -990 -136 -990 1 Dna3
rlabel metal1 -126 -992 -126 -992 1 Aa3
rlabel metal1 -137 -1060 -137 -1060 1 Dna3
rlabel metal1 -107 -1060 -107 -1060 1 Aa3
rlabel metal1 -107 -990 -107 -990 1 Aa3
rlabel metal1 -183 -1266 -183 -1266 1 gnd
rlabel metal1 -153 -1266 -153 -1266 1 gnd
rlabel metal1 -180 -1220 -180 -1220 1 CLK
rlabel metal1 -189 -1103 -189 -1103 1 vdd
rlabel metal1 -150 -1220 -150 -1220 1 CLK
rlabel metal1 -159 -1103 -159 -1103 1 vdd
rlabel metal1 -121 -1197 -121 -1197 1 CLK
rlabel metal1 -128 -1239 -128 -1239 1 gnd
rlabel metal1 -134 -1102 -134 -1102 1 vdd
rlabel metal1 -91 -1197 -91 -1197 1 CLK
rlabel metal1 -98 -1239 -98 -1239 1 gnd
rlabel metal1 -104 -1102 -104 -1102 1 vdd
rlabel metal1 -194 -1162 -194 -1162 1 B3_unlatched
rlabel metal1 -179 -1235 -179 -1235 1 B3_unlatched
rlabel metal1 -191 -1228 -191 -1228 1 Bb3
rlabel metal1 -151 -1235 -151 -1235 1 Bb3
rlabel metal1 -164 -1162 -164 -1162 1 Bb3
rlabel metal1 -133 -1162 -133 -1162 1 Dnb3
rlabel metal1 -123 -1164 -123 -1164 1 Ab3
rlabel metal1 -134 -1232 -134 -1232 1 Dnb3
rlabel metal1 -104 -1232 -104 -1232 1 Ab3
rlabel metal1 -104 -1162 -104 -1162 1 Ab3
rlabel metal1 -191 -213 -191 -213 1 B0_unlatched
rlabel metal1 -219 -1191 -219 -1191 1 gnd
rlabel metal1 -222 -1102 -222 -1102 5 vdd
rlabel metal1 -222 -1019 -222 -1019 1 gnd
rlabel metal1 -225 -930 -225 -930 5 vdd
rlabel metal1 -224 -848 -224 -848 1 gnd
rlabel metal1 -227 -759 -227 -759 5 vdd
rlabel metal1 -227 -677 -227 -677 1 gnd
rlabel metal1 -230 -588 -230 -588 5 vdd
rlabel metal1 -232 -507 -232 -507 1 gnd
rlabel metal1 -235 -418 -235 -418 5 vdd
rlabel metal1 -233 -338 -233 -338 1 gnd
rlabel metal1 -235 -249 -235 -249 1 vdd
rlabel metal1 -234 -80 -234 -80 5 vdd
rlabel metal1 -232 -168 -232 -168 1 gnd
rlabel metal1 -234 3 -234 3 1 gnd
rlabel metal1 -237 92 -237 92 5 vdd
rlabel metal1 -240 35 -240 35 3 Dna0_n
rlabel metal1 -223 35 -223 35 1 Dna0
rlabel metal1 -237 -137 -237 -137 1 Dnb0_n
rlabel metal1 -220 -137 -220 -137 1 Dnb0
rlabel metal1 -238 -306 -238 -306 1 Dna1_n
rlabel metal1 -222 -306 -222 -306 1 Dna1
rlabel metal1 -238 -475 -238 -475 1 Dnb1_n
rlabel metal1 -221 -475 -221 -475 1 Dnb1
rlabel metal1 -233 -645 -233 -645 1 Dna2_n
rlabel metal1 -216 -645 -216 -645 1 Dna2
rlabel metal1 -230 -816 -230 -816 1 Dnb2_n
rlabel metal1 -213 -816 -213 -816 1 Dnb2
rlabel metal1 -228 -987 -228 -987 1 Dna3_n
rlabel metal1 -211 -987 -211 -987 1 Dna3
rlabel metal1 -225 -1159 -225 -1159 1 Dnb3_n
rlabel metal1 -208 -1159 -208 -1159 1 Dnb3
rlabel metal1 -176 -35 -176 -35 1 Dna0_n
rlabel metal1 -173 -206 -173 -206 1 Dnb0_n
rlabel metal1 -175 -375 -175 -375 1 Dna1_n
rlabel metal1 -174 -544 -174 -544 1 Dnb1_n
rlabel metal1 -169 -714 -169 -714 1 Dna2_n
rlabel metal1 -166 -885 -166 -885 1 Dnb2_n
rlabel metal1 -164 -1056 -164 -1056 1 Dna3_n
rlabel metal1 -161 -1228 -161 -1228 1 Dnb3_n
rlabel metal1 -108 29 -108 29 1 A0_n1
rlabel metal1 -105 -142 -105 -142 1 B0_n1
rlabel metal1 -107 -311 -107 -311 1 A1_n1
rlabel metal1 -106 -480 -106 -480 1 B1_n1
rlabel metal1 -101 -650 -101 -650 1 A2_n1
rlabel metal1 -98 -821 -98 -821 1 B2_n1
rlabel metal1 -96 -992 -96 -992 1 A3_n1
rlabel metal1 -93 -1164 -93 -1164 1 B3_n1
rlabel metal1 -90 34 -90 34 1 A0_n1
rlabel metal1 -73 34 -73 34 1 A0
rlabel metal1 -55 34 -55 34 1 B0_n1
rlabel metal1 -39 34 -39 34 1 B0
rlabel metal1 -84 -63 -84 -63 1 A1_n1
rlabel metal1 -70 -63 -70 -63 1 A1
rlabel metal1 -83 -159 -83 -159 1 A2_n1
rlabel metal1 -67 -159 -67 -159 1 A2
rlabel metal1 -78 -256 -78 -256 1 A3_n1
rlabel metal1 -63 -256 -63 -256 1 A3
rlabel metal1 -45 -256 -45 -256 1 B3_n1
rlabel metal1 -29 -256 -29 -256 1 B3
rlabel metal1 -49 -159 -49 -159 1 B2_n1
rlabel metal1 -34 -159 -34 -159 1 B2
rlabel metal1 -50 -63 -50 -63 1 B1_n1
rlabel metal1 -34 -63 -34 -63 1 B1
rlabel metal1 523 1 523 1 1 gnd
rlabel metal1 520 90 520 90 5 vdd
rlabel metal1 523 -170 523 -170 1 gnd
rlabel metal1 520 -81 520 -81 5 vdd
rlabel metal1 524 -339 524 -339 1 gnd
rlabel metal1 521 -250 521 -250 5 vdd
rlabel metal1 524 -507 524 -507 1 gnd
rlabel metal1 521 -418 521 -418 5 vdd
rlabel metal1 525 -678 525 -678 1 gnd
rlabel metal1 522 -589 522 -589 5 vdd
rlabel metal1 553 89 553 89 1 vdd
rlabel metal1 583 89 583 89 1 vdd
rlabel metal1 559 -74 559 -74 1 gnd
rlabel metal1 589 -74 589 -74 1 gnd
rlabel metal1 614 -47 614 -47 1 gnd
rlabel metal1 608 90 608 90 1 vdd
rlabel metal1 644 -47 644 -47 1 gnd
rlabel metal1 638 90 638 90 1 vdd
rlabel metal1 556 -82 556 -82 1 vdd
rlabel metal1 586 -82 586 -82 1 vdd
rlabel metal1 562 -245 562 -245 1 gnd
rlabel metal1 592 -245 592 -245 1 gnd
rlabel metal1 617 -218 617 -218 1 gnd
rlabel metal1 611 -81 611 -81 1 vdd
rlabel metal1 647 -218 647 -218 1 gnd
rlabel metal1 641 -81 641 -81 1 vdd
rlabel metal1 554 -251 554 -251 1 vdd
rlabel metal1 584 -251 584 -251 1 vdd
rlabel metal1 560 -414 560 -414 1 gnd
rlabel metal1 590 -414 590 -414 1 gnd
rlabel metal1 615 -387 615 -387 1 gnd
rlabel metal1 609 -250 609 -250 1 vdd
rlabel metal1 645 -387 645 -387 1 gnd
rlabel metal1 639 -250 639 -250 1 vdd
rlabel metal1 555 -420 555 -420 1 vdd
rlabel metal1 585 -420 585 -420 1 vdd
rlabel metal1 561 -583 561 -583 1 gnd
rlabel metal1 591 -583 591 -583 1 gnd
rlabel metal1 616 -556 616 -556 1 gnd
rlabel metal1 610 -419 610 -419 1 vdd
rlabel metal1 646 -556 646 -556 1 gnd
rlabel metal1 640 -419 640 -419 1 vdd
rlabel metal1 560 -590 560 -590 1 vdd
rlabel metal1 590 -590 590 -590 1 vdd
rlabel metal1 566 -753 566 -753 1 gnd
rlabel metal1 596 -753 596 -753 1 gnd
rlabel metal1 621 -726 621 -726 1 gnd
rlabel metal1 615 -589 615 -589 1 vdd
rlabel metal1 651 -726 651 -726 1 gnd
rlabel metal1 645 -589 645 -589 1 vdd
rlabel metal1 548 30 548 30 1 Sum0_unlatched
rlabel metal1 562 -28 562 -28 1 CLK2
rlabel metal1 551 -36 551 -36 1 Bs0
rlabel metal1 591 -43 591 -43 1 Bs0
rlabel metal1 592 -28 592 -28 1 CLK2
rlabel metal1 578 30 578 30 1 Bs0
rlabel metal1 609 30 609 30 1 Dns0
rlabel metal1 619 28 619 28 1 As0
rlabel metal1 621 -5 621 -5 1 CLK2
rlabel metal1 608 -40 608 -40 1 Dns0
rlabel metal1 638 30 638 30 1 As0
rlabel metal1 638 -40 638 -40 1 As0
rlabel metal1 651 -5 651 -5 1 CLK2
rlabel metal1 563 -43 563 -43 1 Sum0_unlatched
rlabel metal1 551 -141 551 -141 1 Sum1_unlatched
rlabel metal1 565 -199 565 -199 1 CLK2
rlabel metal1 554 -207 554 -207 1 Bs1
rlabel metal1 581 -141 581 -141 1 Bs1
rlabel metal1 594 -214 594 -214 1 Bs1
rlabel metal1 595 -199 595 -199 1 CLK2
rlabel metal1 611 -211 611 -211 1 Dns1
rlabel metal1 624 -176 624 -176 1 CLK2
rlabel metal1 612 -141 612 -141 1 Dns1
rlabel metal1 622 -143 622 -143 1 As1
rlabel metal1 641 -141 641 -141 1 As1
rlabel metal1 641 -211 641 -211 1 As1
rlabel metal1 654 -176 654 -176 1 CLK2
rlabel metal1 566 -214 566 -214 1 Sum1_unlatched
rlabel metal1 549 -310 549 -310 1 Sum2_unlatched
rlabel metal1 564 -383 564 -383 1 Sum2_unlatched
rlabel metal1 563 -368 563 -368 1 CLK2
rlabel metal1 552 -376 552 -376 1 Bs2
rlabel metal1 592 -383 592 -383 1 Bs2
rlabel metal1 593 -368 593 -368 1 CLK2
rlabel metal1 579 -310 579 -310 1 Bs2
rlabel metal1 610 -310 610 -310 1 Dns2
rlabel metal1 622 -345 622 -345 1 CLK2
rlabel metal1 609 -380 609 -380 1 Dns2
rlabel metal1 620 -311 620 -311 1 As2
rlabel metal1 639 -310 639 -310 1 As2
rlabel metal1 639 -380 639 -380 1 As2
rlabel metal1 652 -345 652 -345 1 CLK2
rlabel metal1 550 -479 550 -479 1 Sum3_unlatched
rlabel metal1 564 -537 564 -537 1 CLK2
rlabel metal1 565 -552 565 -552 1 Sum3_unlatched
rlabel metal1 593 -552 593 -552 1 Bs3
rlabel metal1 594 -537 594 -537 1 CLK2
rlabel metal1 610 -549 610 -549 1 Dns3
rlabel metal1 623 -514 623 -514 1 CLK2
rlabel metal1 611 -479 611 -479 1 Dns3
rlabel metal1 621 -481 621 -481 1 As3
rlabel metal1 640 -479 640 -479 1 As3
rlabel metal1 653 -514 653 -514 1 CLK2
rlabel metal1 640 -549 640 -549 1 As3
rlabel metal1 555 -649 555 -649 1 Cout_unlatched
rlabel metal1 570 -722 570 -722 1 Cout_unlatched
rlabel metal1 558 -715 558 -715 1 Bc4
rlabel metal1 569 -707 569 -707 1 CLK2
rlabel metal1 598 -722 598 -722 1 Bc4
rlabel metal1 599 -707 599 -707 1 CLK2
rlabel metal1 615 -719 615 -719 1 Dnc4
rlabel metal1 628 -684 628 -684 1 CLK2
rlabel metal1 616 -649 616 -649 1 Dnc4
rlabel metal1 626 -651 626 -651 1 Ac4
rlabel metal1 645 -649 645 -649 1 Ac4
rlabel metal1 645 -719 645 -719 1 Ac4
rlabel metal1 658 -684 658 -684 1 CLK2
rlabel metal1 580 -479 580 -479 1 Bs3
rlabel metal1 553 -545 553 -545 1 Bs3
rlabel metal1 585 -649 585 -649 1 Bc4
rlabel metal1 517 33 517 33 1 Dns0_n
rlabel metal1 534 33 534 33 1 Dns0
rlabel metal1 581 -36 581 -36 1 Dns0_n
rlabel metal1 517 -138 517 -138 1 Dns1_n
rlabel metal1 534 -138 534 -138 1 Dns1
rlabel metal1 584 -207 584 -207 1 Dns1_n
rlabel metal1 518 -307 518 -307 1 Dns2_n
rlabel metal1 535 -307 535 -307 1 Dns2
rlabel metal1 582 -376 582 -376 1 Dns2_n
rlabel metal1 518 -475 518 -475 1 Dns3_n
rlabel metal1 535 -475 535 -475 1 Dns3
rlabel metal1 583 -545 583 -545 1 Dns3_n
rlabel metal1 519 -646 519 -646 1 Dnc4_n
rlabel metal1 536 -646 536 -646 1 Dnc4
rlabel metal1 588 -715 588 -715 1 Dnc4_n
rlabel metal1 673 1 673 1 1 gnd
rlabel metal1 670 90 670 90 5 vdd
rlabel metal1 676 -170 676 -170 1 gnd
rlabel metal1 673 -81 673 -81 5 vdd
rlabel metal1 674 -339 674 -339 1 gnd
rlabel metal1 671 -250 671 -250 5 vdd
rlabel metal1 675 -508 675 -508 1 gnd
rlabel metal1 672 -419 672 -419 5 vdd
rlabel metal1 680 -678 680 -678 1 gnd
rlabel metal1 677 -589 677 -589 5 vdd
rlabel metal1 684 33 684 33 1 Sum0
rlabel metal1 687 -138 687 -138 1 Sum1
rlabel metal1 685 -307 685 -307 1 Sum2
rlabel metal1 686 -477 686 -477 1 Sum3
rlabel metal1 692 -646 692 -646 7 Cout
<< end >>
