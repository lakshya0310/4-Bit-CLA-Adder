magic
tech scmos
timestamp 1731951454
<< nwell >>
rect -246 1348 -222 1440
rect -246 1237 -222 1329
rect -212 1238 -188 1290
<< ntransistor >>
rect -235 1200 -233 1220
rect -217 1200 -215 1220
rect -201 1209 -199 1229
<< ptransistor >>
rect -235 1354 -233 1434
rect -235 1243 -233 1323
rect -201 1244 -199 1284
<< ndiffusion >>
rect -236 1200 -235 1220
rect -233 1200 -232 1220
rect -218 1200 -217 1220
rect -215 1200 -214 1220
rect -202 1209 -201 1229
rect -199 1209 -198 1229
<< pdiffusion >>
rect -236 1354 -235 1434
rect -233 1354 -232 1434
rect -236 1243 -235 1323
rect -233 1243 -232 1323
rect -202 1244 -201 1284
rect -199 1244 -198 1284
<< ndcontact >>
rect -240 1200 -236 1220
rect -232 1200 -228 1220
rect -222 1200 -218 1220
rect -214 1200 -210 1220
rect -206 1209 -202 1229
rect -198 1209 -194 1229
<< pdcontact >>
rect -240 1354 -236 1434
rect -232 1354 -228 1434
rect -240 1243 -236 1323
rect -232 1243 -228 1323
rect -206 1244 -202 1284
rect -198 1244 -194 1284
<< polysilicon >>
rect -235 1434 -233 1437
rect -235 1341 -233 1354
rect -235 1323 -233 1336
rect -201 1284 -199 1287
rect -235 1233 -233 1243
rect -201 1229 -199 1244
rect -235 1220 -233 1227
rect -217 1220 -215 1227
rect -201 1206 -199 1209
rect -235 1197 -233 1200
rect -217 1197 -215 1200
<< polycontact >>
rect -233 1341 -229 1345
rect -233 1332 -229 1336
rect -205 1232 -201 1236
rect -239 1223 -235 1227
rect -215 1223 -211 1227
<< metal1 >>
rect -246 1438 -222 1442
rect -232 1434 -228 1438
rect -240 1323 -236 1354
rect -229 1341 -227 1345
rect -229 1332 -227 1336
rect -212 1288 -188 1292
rect -206 1284 -202 1288
rect -232 1236 -228 1243
rect -198 1236 -194 1244
rect -232 1232 -205 1236
rect -198 1232 -189 1236
rect -232 1227 -228 1232
rect -198 1229 -194 1232
rect -241 1223 -239 1227
rect -232 1224 -218 1227
rect -232 1220 -228 1224
rect -222 1220 -218 1224
rect -211 1223 -209 1227
rect -206 1204 -202 1209
rect -206 1200 -194 1204
rect -240 1196 -236 1200
rect -214 1196 -210 1200
rect -240 1193 -210 1196
<< labels >>
rlabel metal1 -226 1195 -226 1195 1 gnd
rlabel metal1 -234 1441 -234 1441 5 vdd
rlabel metal1 -202 1202 -202 1202 1 gnd
rlabel metal1 -205 1291 -205 1291 5 vdd
rlabel metal1 -228 1343 -228 1343 1 PC0
rlabel metal1 -228 1334 -228 1334 1 G0
rlabel metal1 -240 1224 -240 1224 1 PC0
rlabel metal1 -210 1225 -210 1225 1 G0
rlabel metal1 -191 1234 -191 1234 7 C1
<< end >>
