magic
tech scmos
timestamp 1731951022
<< nwell >>
rect -463 1276 -439 1328
rect -429 1276 -405 1328
rect -379 1265 -355 1357
rect -349 1265 -325 1357
rect -379 1160 -355 1252
rect -349 1160 -325 1252
<< ntransistor >>
rect -452 1247 -450 1267
rect -418 1247 -416 1267
rect -368 1099 -366 1139
rect -338 1099 -336 1139
rect -368 1044 -366 1084
rect -338 1044 -336 1084
<< ptransistor >>
rect -452 1282 -450 1322
rect -418 1282 -416 1322
rect -368 1271 -366 1351
rect -338 1271 -336 1351
rect -368 1166 -366 1246
rect -338 1166 -336 1246
<< ndiffusion >>
rect -453 1247 -452 1267
rect -450 1247 -449 1267
rect -419 1247 -418 1267
rect -416 1247 -415 1267
rect -369 1099 -368 1139
rect -366 1099 -365 1139
rect -339 1099 -338 1139
rect -336 1099 -335 1139
rect -369 1044 -368 1084
rect -366 1044 -365 1084
rect -339 1044 -338 1084
rect -336 1044 -335 1084
<< pdiffusion >>
rect -453 1282 -452 1322
rect -450 1282 -449 1322
rect -419 1282 -418 1322
rect -416 1282 -415 1322
rect -369 1271 -368 1351
rect -366 1271 -365 1351
rect -339 1271 -338 1351
rect -336 1271 -335 1351
rect -369 1166 -368 1246
rect -366 1166 -365 1246
rect -339 1166 -338 1246
rect -336 1166 -335 1246
<< ndcontact >>
rect -457 1247 -453 1267
rect -449 1247 -445 1267
rect -423 1247 -419 1267
rect -415 1247 -411 1267
rect -373 1099 -369 1139
rect -365 1099 -361 1139
rect -343 1099 -339 1139
rect -335 1099 -331 1139
rect -373 1044 -369 1084
rect -365 1044 -361 1084
rect -343 1044 -339 1084
rect -335 1044 -331 1084
<< pdcontact >>
rect -457 1282 -453 1322
rect -449 1282 -445 1322
rect -423 1282 -419 1322
rect -415 1282 -411 1322
rect -373 1271 -369 1351
rect -365 1271 -361 1351
rect -343 1271 -339 1351
rect -335 1271 -331 1351
rect -373 1166 -369 1246
rect -365 1166 -361 1246
rect -343 1166 -339 1246
rect -335 1166 -331 1246
<< polysilicon >>
rect -368 1351 -366 1354
rect -338 1351 -336 1354
rect -452 1322 -450 1325
rect -418 1322 -416 1325
rect -452 1267 -450 1282
rect -418 1267 -416 1282
rect -368 1260 -366 1271
rect -338 1260 -336 1271
rect -452 1244 -450 1247
rect -418 1244 -416 1247
rect -368 1246 -366 1249
rect -338 1246 -336 1249
rect -368 1155 -366 1166
rect -338 1155 -336 1166
rect -368 1139 -366 1146
rect -338 1139 -336 1146
rect -368 1093 -366 1099
rect -338 1093 -336 1099
rect -368 1084 -366 1087
rect -338 1084 -336 1087
rect -368 1037 -366 1044
rect -338 1037 -336 1044
<< polycontact >>
rect -456 1270 -452 1274
rect -422 1270 -418 1274
rect -372 1260 -368 1264
rect -342 1260 -338 1264
rect -366 1155 -362 1159
rect -336 1155 -332 1159
rect -366 1142 -362 1146
rect -336 1142 -332 1146
rect -366 1037 -362 1041
rect -336 1037 -332 1041
<< metal1 >>
rect -379 1355 -355 1359
rect -349 1355 -325 1359
rect -373 1351 -369 1355
rect -343 1351 -339 1355
rect -463 1326 -439 1330
rect -429 1326 -405 1330
rect -457 1322 -453 1326
rect -423 1322 -419 1326
rect -449 1274 -445 1282
rect -415 1274 -411 1282
rect -460 1270 -456 1274
rect -449 1270 -440 1274
rect -426 1270 -422 1274
rect -415 1270 -407 1274
rect -449 1267 -445 1270
rect -415 1267 -411 1270
rect -374 1260 -372 1264
rect -365 1257 -361 1271
rect -344 1260 -342 1264
rect -335 1257 -331 1271
rect -365 1254 -331 1257
rect -457 1242 -453 1247
rect -423 1242 -419 1247
rect -365 1246 -361 1254
rect -335 1246 -331 1254
rect -457 1238 -445 1242
rect -423 1238 -411 1242
rect -373 1152 -369 1166
rect -362 1155 -360 1159
rect -343 1152 -339 1166
rect -332 1155 -330 1159
rect -373 1149 -339 1152
rect -373 1139 -369 1149
rect -362 1142 -360 1146
rect -343 1139 -339 1149
rect -332 1142 -330 1146
rect -365 1084 -361 1099
rect -335 1084 -331 1099
rect -373 1034 -369 1044
rect -362 1037 -360 1041
rect -343 1034 -339 1044
rect -332 1037 -330 1041
rect -373 1031 -364 1034
rect -343 1031 -334 1034
<< labels >>
rlabel metal1 -453 1240 -453 1240 1 gnd
rlabel metal1 -419 1240 -419 1240 1 gnd
rlabel metal1 -459 1272 -459 1272 1 A0
rlabel metal1 -442 1272 -442 1272 1 A0_n
rlabel metal1 -424 1272 -424 1272 1 B0
rlabel metal1 -408 1272 -408 1272 1 B0_n
rlabel metal1 -456 1329 -456 1329 5 vdd
rlabel metal1 -422 1329 -422 1329 5 vdd
rlabel metal1 -372 1358 -372 1358 5 vdd
rlabel metal1 -343 1358 -343 1358 5 vdd
rlabel metal1 -370 1033 -370 1033 1 gnd
rlabel metal1 -340 1033 -340 1033 1 gnd
rlabel metal1 -373 1262 -373 1262 1 A0
rlabel metal1 -343 1262 -343 1262 1 B0
rlabel metal1 -361 1157 -361 1157 1 A0_n
rlabel metal1 -331 1157 -331 1157 1 B0_n
rlabel metal1 -361 1144 -361 1144 1 A0
rlabel metal1 -331 1144 -331 1144 1 A0_n
rlabel metal1 -361 1039 -361 1039 1 B0
rlabel metal1 -331 1039 -331 1039 1 B0_n
rlabel metal1 -341 1151 -341 1151 1 P0
<< end >>
