magic
tech scmos
timestamp 1731951280
<< nwell >>
rect -286 1406 -262 1458
rect -256 1406 -232 1458
rect -226 1406 -202 1458
<< ntransistor >>
rect -275 1349 -273 1389
rect -215 1377 -213 1397
rect -275 1298 -273 1338
<< ptransistor >>
rect -275 1412 -273 1452
rect -245 1412 -243 1452
rect -215 1412 -213 1452
<< ndiffusion >>
rect -276 1349 -275 1389
rect -273 1349 -272 1389
rect -216 1377 -215 1397
rect -213 1377 -212 1397
rect -276 1298 -275 1338
rect -273 1298 -272 1338
<< pdiffusion >>
rect -276 1412 -275 1452
rect -273 1412 -272 1452
rect -246 1412 -245 1452
rect -243 1412 -242 1452
rect -216 1412 -215 1452
rect -213 1412 -212 1452
<< ndcontact >>
rect -280 1349 -276 1389
rect -272 1349 -268 1389
rect -220 1377 -216 1397
rect -212 1377 -208 1397
rect -280 1298 -276 1338
rect -272 1298 -268 1338
<< pdcontact >>
rect -280 1412 -276 1452
rect -272 1412 -268 1452
rect -250 1412 -246 1452
rect -242 1412 -238 1452
rect -220 1412 -216 1452
rect -212 1412 -208 1452
<< polysilicon >>
rect -275 1452 -273 1455
rect -245 1452 -243 1455
rect -215 1452 -213 1455
rect -275 1401 -273 1412
rect -245 1401 -243 1412
rect -215 1397 -213 1412
rect -275 1389 -273 1396
rect -215 1374 -213 1377
rect -275 1346 -273 1349
rect -275 1338 -273 1341
rect -275 1291 -273 1298
<< polycontact >>
rect -279 1401 -275 1405
rect -249 1401 -245 1405
rect -219 1400 -215 1404
rect -279 1392 -275 1396
rect -279 1291 -275 1295
<< metal1 >>
rect -286 1456 -232 1460
rect -226 1456 -202 1460
rect -280 1452 -276 1456
rect -250 1452 -246 1456
rect -220 1452 -216 1456
rect -281 1401 -279 1405
rect -272 1398 -268 1412
rect -251 1401 -249 1405
rect -242 1404 -238 1412
rect -212 1404 -208 1412
rect -242 1400 -219 1404
rect -212 1400 -203 1404
rect -242 1398 -238 1400
rect -281 1392 -279 1396
rect -272 1395 -238 1398
rect -212 1397 -208 1400
rect -272 1389 -268 1395
rect -220 1372 -216 1377
rect -220 1368 -208 1372
rect -280 1338 -276 1349
rect -281 1291 -279 1295
rect -272 1288 -268 1298
rect -281 1285 -268 1288
<< labels >>
rlabel metal1 -273 1287 -273 1287 1 gnd
rlabel metal1 -216 1370 -216 1370 1 gnd
rlabel metal1 -219 1459 -219 1459 5 vdd
rlabel metal1 -261 1459 -261 1459 5 vdd
rlabel metal1 -280 1403 -280 1403 1 A0
rlabel metal1 -250 1403 -250 1403 1 B0
rlabel metal1 -280 1394 -280 1394 1 A0
rlabel metal1 -280 1293 -280 1293 1 B0
rlabel nwell -204 1411 -204 1411 1 G0
<< end >>
