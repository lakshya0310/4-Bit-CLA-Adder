magic
tech scmos
timestamp 1732001842
<< nwell >>
rect 1963 2249 1987 2301
rect 1993 2245 2017 2300
rect 2023 2245 2047 2300
rect 2053 2245 2077 2300
rect 2083 2245 2107 2300
rect 2113 2249 2137 2301
rect 1993 2187 2017 2239
rect 2023 2187 2047 2239
<< ntransistor >>
rect 1974 2220 1976 2240
rect 2064 2213 2066 2233
rect 2094 2213 2096 2233
rect 2124 2220 2126 2240
rect 2064 2178 2066 2198
rect 2094 2178 2096 2198
rect 2004 2144 2006 2164
rect 2034 2144 2036 2164
<< ptransistor >>
rect 1974 2255 1976 2295
rect 2004 2254 2006 2294
rect 2034 2254 2036 2294
rect 2064 2254 2066 2294
rect 2094 2254 2096 2294
rect 2124 2255 2126 2295
rect 2004 2193 2006 2233
rect 2034 2193 2036 2233
<< ndiffusion >>
rect 1973 2220 1974 2240
rect 1976 2220 1977 2240
rect 2063 2213 2064 2233
rect 2066 2213 2067 2233
rect 2093 2213 2094 2233
rect 2096 2213 2097 2233
rect 2123 2220 2124 2240
rect 2126 2220 2127 2240
rect 2063 2178 2064 2198
rect 2066 2178 2067 2198
rect 2093 2178 2094 2198
rect 2096 2178 2097 2198
rect 2003 2144 2004 2164
rect 2006 2144 2007 2164
rect 2033 2144 2034 2164
rect 2036 2144 2037 2164
<< pdiffusion >>
rect 1973 2255 1974 2295
rect 1976 2255 1977 2295
rect 2003 2254 2004 2294
rect 2006 2254 2007 2294
rect 2033 2254 2034 2294
rect 2036 2254 2037 2294
rect 2063 2254 2064 2294
rect 2066 2254 2067 2294
rect 2093 2254 2094 2294
rect 2096 2254 2097 2294
rect 2123 2255 2124 2295
rect 2126 2255 2127 2295
rect 2003 2193 2004 2233
rect 2006 2193 2007 2233
rect 2033 2193 2034 2233
rect 2036 2193 2037 2233
<< ndcontact >>
rect 1969 2220 1973 2240
rect 1977 2220 1981 2240
rect 2059 2213 2063 2233
rect 2067 2213 2071 2233
rect 2089 2213 2093 2233
rect 2097 2213 2101 2233
rect 2119 2220 2123 2240
rect 2127 2220 2131 2240
rect 2059 2178 2063 2198
rect 2067 2178 2071 2198
rect 2089 2178 2093 2198
rect 2097 2178 2101 2198
rect 1999 2144 2003 2164
rect 2007 2144 2011 2164
rect 2029 2144 2033 2164
rect 2037 2144 2041 2164
<< pdcontact >>
rect 1969 2255 1973 2295
rect 1977 2255 1981 2295
rect 1999 2254 2003 2294
rect 2007 2254 2011 2294
rect 2029 2254 2033 2294
rect 2037 2254 2041 2294
rect 2059 2254 2063 2294
rect 2067 2254 2071 2294
rect 2089 2254 2093 2294
rect 2097 2254 2101 2294
rect 2119 2255 2123 2295
rect 2127 2255 2131 2295
rect 1999 2193 2003 2233
rect 2007 2193 2011 2233
rect 2029 2193 2033 2233
rect 2037 2193 2041 2233
<< polysilicon >>
rect 1974 2295 1976 2298
rect 2004 2294 2006 2297
rect 2034 2294 2036 2297
rect 2064 2294 2066 2297
rect 2094 2294 2096 2297
rect 2124 2295 2126 2298
rect 1974 2240 1976 2255
rect 2004 2240 2006 2254
rect 2034 2240 2036 2254
rect 2064 2240 2066 2254
rect 2094 2240 2096 2254
rect 2124 2240 2126 2255
rect 2004 2233 2006 2236
rect 2034 2233 2036 2236
rect 2064 2233 2066 2236
rect 2094 2233 2096 2236
rect 1974 2217 1976 2220
rect 2124 2217 2126 2220
rect 2064 2205 2066 2213
rect 2094 2205 2096 2213
rect 2064 2198 2066 2201
rect 2094 2198 2096 2201
rect 2004 2182 2006 2193
rect 2034 2182 2036 2193
rect 2004 2164 2006 2171
rect 2034 2164 2036 2171
rect 2064 2170 2066 2178
rect 2094 2170 2096 2178
rect 2004 2141 2006 2144
rect 2034 2141 2036 2144
<< polycontact >>
rect 1970 2243 1974 2247
rect 2000 2240 2004 2244
rect 2030 2240 2034 2244
rect 2060 2240 2064 2244
rect 2090 2240 2094 2244
rect 2120 2243 2124 2247
rect 2066 2205 2070 2209
rect 2096 2205 2100 2209
rect 2006 2182 2010 2186
rect 2036 2182 2040 2186
rect 2006 2167 2010 2171
rect 2036 2167 2040 2171
rect 2060 2170 2064 2174
rect 2090 2170 2094 2174
<< metal1 >>
rect 1963 2299 1987 2303
rect 1993 2300 2017 2303
rect 2023 2300 2047 2303
rect 2053 2300 2077 2303
rect 2083 2300 2107 2303
rect 1969 2295 1973 2299
rect 1977 2247 1981 2255
rect 1999 2294 2003 2300
rect 2029 2294 2033 2300
rect 2059 2294 2063 2300
rect 2089 2294 2093 2300
rect 2113 2299 2137 2303
rect 2119 2295 2123 2299
rect 1966 2243 1970 2247
rect 1977 2243 1986 2247
rect 1977 2240 1981 2243
rect 1997 2240 2000 2244
rect 2007 2233 2011 2254
rect 2027 2240 2030 2244
rect 2037 2233 2041 2254
rect 2057 2240 2060 2244
rect 2067 2233 2071 2254
rect 2087 2240 2090 2244
rect 2097 2243 2101 2254
rect 2127 2247 2131 2255
rect 2113 2243 2120 2247
rect 2127 2243 2136 2247
rect 2097 2239 2116 2243
rect 2127 2240 2131 2243
rect 2097 2233 2101 2239
rect 1969 2215 1973 2220
rect 1969 2211 1981 2215
rect 2119 2215 2123 2220
rect 2059 2198 2063 2213
rect 2070 2205 2073 2209
rect 2089 2198 2093 2213
rect 2119 2211 2131 2215
rect 2100 2205 2103 2209
rect 1999 2164 2003 2193
rect 2010 2182 2014 2186
rect 2010 2167 2014 2171
rect 2029 2164 2033 2193
rect 2040 2182 2044 2186
rect 2040 2167 2046 2171
rect 2057 2170 2060 2174
rect 2067 2167 2071 2178
rect 2087 2170 2090 2174
rect 2097 2167 2101 2178
rect 2057 2164 2071 2167
rect 2087 2164 2101 2167
rect 2007 2140 2011 2144
rect 2037 2140 2041 2144
rect 1999 2137 2011 2140
rect 2029 2137 2041 2140
<< labels >>
rlabel metal1 1973 2213 1973 2213 1 gnd
rlabel metal1 1970 2302 1970 2302 5 vdd
rlabel metal1 2003 2301 2003 2301 1 vdd
rlabel metal1 2033 2301 2033 2301 1 vdd
rlabel metal1 2009 2138 2009 2138 1 gnd
rlabel metal1 2039 2138 2039 2138 1 gnd
rlabel metal1 2064 2165 2064 2165 1 gnd
rlabel metal1 2058 2302 2058 2302 1 vdd
rlabel metal1 2094 2165 2094 2165 1 gnd
rlabel metal1 2088 2302 2088 2302 1 vdd
rlabel metal1 1998 2242 1998 2242 1 Sum0_unlatched
rlabel metal1 2012 2184 2012 2184 1 CLK2
rlabel metal1 2001 2176 2001 2176 1 Bs0
rlabel metal1 2041 2169 2041 2169 1 Bs0
rlabel metal1 2042 2184 2042 2184 1 CLK2
rlabel metal1 2028 2242 2028 2242 1 Bs0
rlabel metal1 2059 2242 2059 2242 1 Dns0
rlabel metal1 2069 2240 2069 2240 1 As0
rlabel metal1 2071 2207 2071 2207 1 CLK2
rlabel metal1 2058 2172 2058 2172 1 Dns0
rlabel metal1 2088 2242 2088 2242 1 As0
rlabel metal1 2088 2172 2088 2172 1 As0
rlabel metal1 2101 2207 2101 2207 1 CLK2
rlabel metal1 2013 2169 2013 2169 1 Sum0_unlatched
rlabel metal1 1967 2245 1967 2245 1 Dns0_n
rlabel metal1 1984 2245 1984 2245 1 Dns0
rlabel metal1 2031 2176 2031 2176 1 Dns0_n
rlabel metal1 2123 2213 2123 2213 1 gnd
rlabel metal1 2120 2302 2120 2302 5 vdd
rlabel metal1 2134 2245 2134 2245 1 Sum0
<< end >>
